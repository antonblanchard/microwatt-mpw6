VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM512
  CLASS BLOCK ;
  FOREIGN RAM512 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1583.780 BY 987.360 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 520.920 1583.780 521.520 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 575.320 1583.780 575.920 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 630.400 1583.780 631.000 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 685.480 1583.780 686.080 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 739.880 1583.780 740.480 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 794.960 1583.780 795.560 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 850.040 1583.780 850.640 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 904.440 1583.780 905.040 ;
    END
  END A0[7]
  PIN A0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 959.520 1583.780 960.120 ;
    END
  END A0[8]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 2.000 494.320 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 0.000 556.510 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 0.000 655.410 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 0.000 705.090 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 0.000 779.150 2.000 ;
    END
  END Di0[31]
  PIN Di0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 0.000 803.990 2.000 ;
    END
  END Di0[32]
  PIN Di0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 0.000 828.830 2.000 ;
    END
  END Di0[33]
  PIN Di0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 2.000 ;
    END
  END Di0[34]
  PIN Di0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 0.000 878.050 2.000 ;
    END
  END Di0[35]
  PIN Di0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 0.000 902.890 2.000 ;
    END
  END Di0[36]
  PIN Di0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 2.000 ;
    END
  END Di0[37]
  PIN Di0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 0.000 952.570 2.000 ;
    END
  END Di0[38]
  PIN Di0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 0.000 977.410 2.000 ;
    END
  END Di0[39]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 2.000 ;
    END
  END Di0[3]
  PIN Di0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 0.000 1001.790 2.000 ;
    END
  END Di0[40]
  PIN Di0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 0.000 1026.630 2.000 ;
    END
  END Di0[41]
  PIN Di0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 0.000 1051.470 2.000 ;
    END
  END Di0[42]
  PIN Di0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.030 0.000 1076.310 2.000 ;
    END
  END Di0[43]
  PIN Di0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.870 0.000 1101.150 2.000 ;
    END
  END Di0[44]
  PIN Di0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.250 0.000 1125.530 2.000 ;
    END
  END Di0[45]
  PIN Di0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 0.000 1150.370 2.000 ;
    END
  END Di0[46]
  PIN Di0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.930 0.000 1175.210 2.000 ;
    END
  END Di0[47]
  PIN Di0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.770 0.000 1200.050 2.000 ;
    END
  END Di0[48]
  PIN Di0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.610 0.000 1224.890 2.000 ;
    END
  END Di0[49]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 2.000 ;
    END
  END Di0[4]
  PIN Di0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.990 0.000 1249.270 2.000 ;
    END
  END Di0[50]
  PIN Di0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 0.000 1274.110 2.000 ;
    END
  END Di0[51]
  PIN Di0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.670 0.000 1298.950 2.000 ;
    END
  END Di0[52]
  PIN Di0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 2.000 ;
    END
  END Di0[53]
  PIN Di0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.350 0.000 1348.630 2.000 ;
    END
  END Di0[54]
  PIN Di0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.730 0.000 1373.010 2.000 ;
    END
  END Di0[55]
  PIN Di0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 0.000 1397.850 2.000 ;
    END
  END Di0[56]
  PIN Di0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.410 0.000 1422.690 2.000 ;
    END
  END Di0[57]
  PIN Di0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.250 0.000 1447.530 2.000 ;
    END
  END Di0[58]
  PIN Di0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.090 0.000 1472.370 2.000 ;
    END
  END Di0[59]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 2.000 ;
    END
  END Di0[5]
  PIN Di0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.470 0.000 1496.750 2.000 ;
    END
  END Di0[60]
  PIN Di0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.310 0.000 1521.590 2.000 ;
    END
  END Di0[61]
  PIN Di0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.150 0.000 1546.430 2.000 ;
    END
  END Di0[62]
  PIN Di0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.990 0.000 1571.270 2.000 ;
    END
  END Di0[63]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 985.360 12.330 987.360 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 985.360 259.350 987.360 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 985.360 284.190 987.360 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 985.360 309.030 987.360 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 985.360 333.870 987.360 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 985.360 358.710 987.360 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 985.360 383.090 987.360 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 985.360 407.930 987.360 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 985.360 432.770 987.360 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 985.360 457.610 987.360 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 985.360 482.450 987.360 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 985.360 36.710 987.360 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 985.360 506.830 987.360 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 985.360 531.670 987.360 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 985.360 556.510 987.360 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 985.360 581.350 987.360 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 985.360 606.190 987.360 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 985.360 630.570 987.360 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 985.360 655.410 987.360 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 985.360 680.250 987.360 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 985.360 705.090 987.360 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 985.360 729.930 987.360 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 985.360 61.550 987.360 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 985.360 754.310 987.360 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 985.360 779.150 987.360 ;
    END
  END Do0[31]
  PIN Do0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 985.360 803.990 987.360 ;
    END
  END Do0[32]
  PIN Do0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 985.360 828.830 987.360 ;
    END
  END Do0[33]
  PIN Do0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 985.360 853.670 987.360 ;
    END
  END Do0[34]
  PIN Do0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 985.360 878.050 987.360 ;
    END
  END Do0[35]
  PIN Do0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 985.360 902.890 987.360 ;
    END
  END Do0[36]
  PIN Do0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 985.360 927.730 987.360 ;
    END
  END Do0[37]
  PIN Do0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 985.360 952.570 987.360 ;
    END
  END Do0[38]
  PIN Do0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 985.360 977.410 987.360 ;
    END
  END Do0[39]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 985.360 86.390 987.360 ;
    END
  END Do0[3]
  PIN Do0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 985.360 1001.790 987.360 ;
    END
  END Do0[40]
  PIN Do0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 985.360 1026.630 987.360 ;
    END
  END Do0[41]
  PIN Do0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 985.360 1051.470 987.360 ;
    END
  END Do0[42]
  PIN Do0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.030 985.360 1076.310 987.360 ;
    END
  END Do0[43]
  PIN Do0[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.870 985.360 1101.150 987.360 ;
    END
  END Do0[44]
  PIN Do0[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.250 985.360 1125.530 987.360 ;
    END
  END Do0[45]
  PIN Do0[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 985.360 1150.370 987.360 ;
    END
  END Do0[46]
  PIN Do0[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.930 985.360 1175.210 987.360 ;
    END
  END Do0[47]
  PIN Do0[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.770 985.360 1200.050 987.360 ;
    END
  END Do0[48]
  PIN Do0[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.610 985.360 1224.890 987.360 ;
    END
  END Do0[49]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 985.360 111.230 987.360 ;
    END
  END Do0[4]
  PIN Do0[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.990 985.360 1249.270 987.360 ;
    END
  END Do0[50]
  PIN Do0[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 985.360 1274.110 987.360 ;
    END
  END Do0[51]
  PIN Do0[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.670 985.360 1298.950 987.360 ;
    END
  END Do0[52]
  PIN Do0[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 985.360 1323.790 987.360 ;
    END
  END Do0[53]
  PIN Do0[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.350 985.360 1348.630 987.360 ;
    END
  END Do0[54]
  PIN Do0[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.730 985.360 1373.010 987.360 ;
    END
  END Do0[55]
  PIN Do0[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 985.360 1397.850 987.360 ;
    END
  END Do0[56]
  PIN Do0[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.410 985.360 1422.690 987.360 ;
    END
  END Do0[57]
  PIN Do0[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.250 985.360 1447.530 987.360 ;
    END
  END Do0[58]
  PIN Do0[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.090 985.360 1472.370 987.360 ;
    END
  END Do0[59]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 985.360 135.610 987.360 ;
    END
  END Do0[5]
  PIN Do0[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.470 985.360 1496.750 987.360 ;
    END
  END Do0[60]
  PIN Do0[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.310 985.360 1521.590 987.360 ;
    END
  END Do0[61]
  PIN Do0[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.150 985.360 1546.430 987.360 ;
    END
  END Do0[62]
  PIN Do0[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.990 985.360 1571.270 987.360 ;
    END
  END Do0[63]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 985.360 160.450 987.360 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 985.360 185.290 987.360 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 985.360 210.130 987.360 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 985.360 234.970 987.360 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 27.240 1583.780 27.840 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 113.690 100.400 116.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 293.690 100.400 296.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 473.690 100.400 476.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.690 100.400 656.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 833.690 100.400 836.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.690 100.400 1016.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1193.690 100.400 1196.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1373.690 100.400 1376.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1553.690 100.400 1556.790 886.960 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.690 100.400 26.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.690 100.400 206.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 383.690 100.400 386.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 563.690 100.400 566.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 743.690 100.400 746.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 923.690 100.400 926.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1103.690 100.400 1106.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.690 100.400 1286.790 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 1463.690 100.400 1466.790 886.960 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 81.640 1583.780 82.240 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 136.720 1583.780 137.320 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 191.800 1583.780 192.400 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 246.200 1583.780 246.800 ;
    END
  END WE0[3]
  PIN WE0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 301.280 1583.780 301.880 ;
    END
  END WE0[4]
  PIN WE0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 356.360 1583.780 356.960 ;
    END
  END WE0[5]
  PIN WE0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 410.760 1583.780 411.360 ;
    END
  END WE0[6]
  PIN WE0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1581.780 465.840 1583.780 466.440 ;
    END
  END WE0[7]
  OBS
      LAYER li1 ;
        RECT 20.240 100.555 1563.540 886.805 ;
      LAYER met1 ;
        RECT 1.450 0.380 1580.950 987.320 ;
      LAYER met2 ;
        RECT 1.480 985.080 11.770 987.350 ;
        RECT 12.610 985.080 36.150 987.350 ;
        RECT 36.990 985.080 60.990 987.350 ;
        RECT 61.830 985.080 85.830 987.350 ;
        RECT 86.670 985.080 110.670 987.350 ;
        RECT 111.510 985.080 135.050 987.350 ;
        RECT 135.890 985.080 159.890 987.350 ;
        RECT 160.730 985.080 184.730 987.350 ;
        RECT 185.570 985.080 209.570 987.350 ;
        RECT 210.410 985.080 234.410 987.350 ;
        RECT 235.250 985.080 258.790 987.350 ;
        RECT 259.630 985.080 283.630 987.350 ;
        RECT 284.470 985.080 308.470 987.350 ;
        RECT 309.310 985.080 333.310 987.350 ;
        RECT 334.150 985.080 358.150 987.350 ;
        RECT 358.990 985.080 382.530 987.350 ;
        RECT 383.370 985.080 407.370 987.350 ;
        RECT 408.210 985.080 432.210 987.350 ;
        RECT 433.050 985.080 457.050 987.350 ;
        RECT 457.890 985.080 481.890 987.350 ;
        RECT 482.730 985.080 506.270 987.350 ;
        RECT 507.110 985.080 531.110 987.350 ;
        RECT 531.950 985.080 555.950 987.350 ;
        RECT 556.790 985.080 580.790 987.350 ;
        RECT 581.630 985.080 605.630 987.350 ;
        RECT 606.470 985.080 630.010 987.350 ;
        RECT 630.850 985.080 654.850 987.350 ;
        RECT 655.690 985.080 679.690 987.350 ;
        RECT 680.530 985.080 704.530 987.350 ;
        RECT 705.370 985.080 729.370 987.350 ;
        RECT 730.210 985.080 753.750 987.350 ;
        RECT 754.590 985.080 778.590 987.350 ;
        RECT 779.430 985.080 803.430 987.350 ;
        RECT 804.270 985.080 828.270 987.350 ;
        RECT 829.110 985.080 853.110 987.350 ;
        RECT 853.950 985.080 877.490 987.350 ;
        RECT 878.330 985.080 902.330 987.350 ;
        RECT 903.170 985.080 927.170 987.350 ;
        RECT 928.010 985.080 952.010 987.350 ;
        RECT 952.850 985.080 976.850 987.350 ;
        RECT 977.690 985.080 1001.230 987.350 ;
        RECT 1002.070 985.080 1026.070 987.350 ;
        RECT 1026.910 985.080 1050.910 987.350 ;
        RECT 1051.750 985.080 1075.750 987.350 ;
        RECT 1076.590 985.080 1100.590 987.350 ;
        RECT 1101.430 985.080 1124.970 987.350 ;
        RECT 1125.810 985.080 1149.810 987.350 ;
        RECT 1150.650 985.080 1174.650 987.350 ;
        RECT 1175.490 985.080 1199.490 987.350 ;
        RECT 1200.330 985.080 1224.330 987.350 ;
        RECT 1225.170 985.080 1248.710 987.350 ;
        RECT 1249.550 985.080 1273.550 987.350 ;
        RECT 1274.390 985.080 1298.390 987.350 ;
        RECT 1299.230 985.080 1323.230 987.350 ;
        RECT 1324.070 985.080 1348.070 987.350 ;
        RECT 1348.910 985.080 1372.450 987.350 ;
        RECT 1373.290 985.080 1397.290 987.350 ;
        RECT 1398.130 985.080 1422.130 987.350 ;
        RECT 1422.970 985.080 1446.970 987.350 ;
        RECT 1447.810 985.080 1471.810 987.350 ;
        RECT 1472.650 985.080 1496.190 987.350 ;
        RECT 1497.030 985.080 1521.030 987.350 ;
        RECT 1521.870 985.080 1545.870 987.350 ;
        RECT 1546.710 985.080 1570.710 987.350 ;
        RECT 1571.550 985.080 1580.920 987.350 ;
        RECT 1.480 2.280 1580.920 985.080 ;
        RECT 1.480 0.155 11.770 2.280 ;
        RECT 12.610 0.155 36.150 2.280 ;
        RECT 36.990 0.155 60.990 2.280 ;
        RECT 61.830 0.155 85.830 2.280 ;
        RECT 86.670 0.155 110.670 2.280 ;
        RECT 111.510 0.155 135.050 2.280 ;
        RECT 135.890 0.155 159.890 2.280 ;
        RECT 160.730 0.155 184.730 2.280 ;
        RECT 185.570 0.155 209.570 2.280 ;
        RECT 210.410 0.155 234.410 2.280 ;
        RECT 235.250 0.155 258.790 2.280 ;
        RECT 259.630 0.155 283.630 2.280 ;
        RECT 284.470 0.155 308.470 2.280 ;
        RECT 309.310 0.155 333.310 2.280 ;
        RECT 334.150 0.155 358.150 2.280 ;
        RECT 358.990 0.155 382.530 2.280 ;
        RECT 383.370 0.155 407.370 2.280 ;
        RECT 408.210 0.155 432.210 2.280 ;
        RECT 433.050 0.155 457.050 2.280 ;
        RECT 457.890 0.155 481.890 2.280 ;
        RECT 482.730 0.155 506.270 2.280 ;
        RECT 507.110 0.155 531.110 2.280 ;
        RECT 531.950 0.155 555.950 2.280 ;
        RECT 556.790 0.155 580.790 2.280 ;
        RECT 581.630 0.155 605.630 2.280 ;
        RECT 606.470 0.155 630.010 2.280 ;
        RECT 630.850 0.155 654.850 2.280 ;
        RECT 655.690 0.155 679.690 2.280 ;
        RECT 680.530 0.155 704.530 2.280 ;
        RECT 705.370 0.155 729.370 2.280 ;
        RECT 730.210 0.155 753.750 2.280 ;
        RECT 754.590 0.155 778.590 2.280 ;
        RECT 779.430 0.155 803.430 2.280 ;
        RECT 804.270 0.155 828.270 2.280 ;
        RECT 829.110 0.155 853.110 2.280 ;
        RECT 853.950 0.155 877.490 2.280 ;
        RECT 878.330 0.155 902.330 2.280 ;
        RECT 903.170 0.155 927.170 2.280 ;
        RECT 928.010 0.155 952.010 2.280 ;
        RECT 952.850 0.155 976.850 2.280 ;
        RECT 977.690 0.155 1001.230 2.280 ;
        RECT 1002.070 0.155 1026.070 2.280 ;
        RECT 1026.910 0.155 1050.910 2.280 ;
        RECT 1051.750 0.155 1075.750 2.280 ;
        RECT 1076.590 0.155 1100.590 2.280 ;
        RECT 1101.430 0.155 1124.970 2.280 ;
        RECT 1125.810 0.155 1149.810 2.280 ;
        RECT 1150.650 0.155 1174.650 2.280 ;
        RECT 1175.490 0.155 1199.490 2.280 ;
        RECT 1200.330 0.155 1224.330 2.280 ;
        RECT 1225.170 0.155 1248.710 2.280 ;
        RECT 1249.550 0.155 1273.550 2.280 ;
        RECT 1274.390 0.155 1298.390 2.280 ;
        RECT 1299.230 0.155 1323.230 2.280 ;
        RECT 1324.070 0.155 1348.070 2.280 ;
        RECT 1348.910 0.155 1372.450 2.280 ;
        RECT 1373.290 0.155 1397.290 2.280 ;
        RECT 1398.130 0.155 1422.130 2.280 ;
        RECT 1422.970 0.155 1446.970 2.280 ;
        RECT 1447.810 0.155 1471.810 2.280 ;
        RECT 1472.650 0.155 1496.190 2.280 ;
        RECT 1497.030 0.155 1521.030 2.280 ;
        RECT 1521.870 0.155 1545.870 2.280 ;
        RECT 1546.710 0.155 1570.710 2.280 ;
        RECT 1571.550 0.155 1580.920 2.280 ;
      LAYER met3 ;
        RECT 1.905 960.520 1581.780 987.185 ;
        RECT 1.905 959.120 1581.380 960.520 ;
        RECT 1.905 905.440 1581.780 959.120 ;
        RECT 1.905 904.040 1581.380 905.440 ;
        RECT 1.905 851.040 1581.780 904.040 ;
        RECT 1.905 849.640 1581.380 851.040 ;
        RECT 1.905 795.960 1581.780 849.640 ;
        RECT 1.905 794.560 1581.380 795.960 ;
        RECT 1.905 740.880 1581.780 794.560 ;
        RECT 1.905 739.480 1581.380 740.880 ;
        RECT 1.905 686.480 1581.780 739.480 ;
        RECT 1.905 685.080 1581.380 686.480 ;
        RECT 1.905 631.400 1581.780 685.080 ;
        RECT 1.905 630.000 1581.380 631.400 ;
        RECT 1.905 576.320 1581.780 630.000 ;
        RECT 1.905 574.920 1581.380 576.320 ;
        RECT 1.905 521.920 1581.780 574.920 ;
        RECT 1.905 520.520 1581.380 521.920 ;
        RECT 1.905 494.720 1581.780 520.520 ;
        RECT 2.400 493.320 1581.780 494.720 ;
        RECT 1.905 466.840 1581.780 493.320 ;
        RECT 1.905 465.440 1581.380 466.840 ;
        RECT 1.905 411.760 1581.780 465.440 ;
        RECT 1.905 410.360 1581.380 411.760 ;
        RECT 1.905 357.360 1581.780 410.360 ;
        RECT 1.905 355.960 1581.380 357.360 ;
        RECT 1.905 302.280 1581.780 355.960 ;
        RECT 1.905 300.880 1581.380 302.280 ;
        RECT 1.905 247.200 1581.780 300.880 ;
        RECT 1.905 245.800 1581.380 247.200 ;
        RECT 1.905 192.800 1581.780 245.800 ;
        RECT 1.905 191.400 1581.380 192.800 ;
        RECT 1.905 137.720 1581.780 191.400 ;
        RECT 1.905 136.320 1581.380 137.720 ;
        RECT 1.905 82.640 1581.780 136.320 ;
        RECT 1.905 81.240 1581.380 82.640 ;
        RECT 1.905 28.240 1581.780 81.240 ;
        RECT 1.905 26.840 1581.380 28.240 ;
        RECT 1.905 0.175 1581.780 26.840 ;
      LAYER met4 ;
        RECT 13.175 887.360 1569.225 987.185 ;
        RECT 13.175 100.000 23.290 887.360 ;
        RECT 27.190 100.000 113.290 887.360 ;
        RECT 117.190 100.000 203.290 887.360 ;
        RECT 207.190 100.000 293.290 887.360 ;
        RECT 297.190 100.000 383.290 887.360 ;
        RECT 387.190 100.000 473.290 887.360 ;
        RECT 477.190 100.000 563.290 887.360 ;
        RECT 567.190 100.000 653.290 887.360 ;
        RECT 657.190 100.000 743.290 887.360 ;
        RECT 747.190 100.000 833.290 887.360 ;
        RECT 837.190 100.000 923.290 887.360 ;
        RECT 927.190 100.000 1013.290 887.360 ;
        RECT 1017.190 100.000 1103.290 887.360 ;
        RECT 1107.190 100.000 1193.290 887.360 ;
        RECT 1197.190 100.000 1283.290 887.360 ;
        RECT 1287.190 100.000 1373.290 887.360 ;
        RECT 1377.190 100.000 1463.290 887.360 ;
        RECT 1467.190 100.000 1553.290 887.360 ;
        RECT 1557.190 100.000 1569.225 887.360 ;
        RECT 13.175 0.855 1569.225 100.000 ;
  END
END RAM512
END LIBRARY

