* NGSPICE file created from multiply_add_64x64.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fa_2 abstract view
.subckt sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fa_1 abstract view
.subckt sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_1 abstract view
.subckt sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_2 abstract view
.subckt sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_4 abstract view
.subckt sky130_fd_sc_hd__ha_4 A B VGND VNB VPB VPWR COUT SUM
.ends

.subckt multiply_add_64x64 VGND VPWR a[0] a[10] a[11] a[12] a[13] a[14] a[15] a[16]
+ a[17] a[18] a[19] a[1] a[20] a[21] a[22] a[23] a[24] a[25] a[26] a[27] a[28] a[29]
+ a[2] a[30] a[31] a[32] a[33] a[34] a[35] a[36] a[37] a[38] a[39] a[3] a[40] a[41]
+ a[42] a[43] a[44] a[45] a[46] a[47] a[48] a[49] a[4] a[50] a[51] a[52] a[53] a[54]
+ a[55] a[56] a[57] a[58] a[59] a[5] a[60] a[61] a[62] a[63] a[6] a[7] a[8] a[9] b[0]
+ b[10] b[11] b[12] b[13] b[14] b[15] b[16] b[17] b[18] b[19] b[1] b[20] b[21] b[22]
+ b[23] b[24] b[25] b[26] b[27] b[28] b[29] b[2] b[30] b[31] b[32] b[33] b[34] b[35]
+ b[36] b[37] b[38] b[39] b[3] b[40] b[41] b[42] b[43] b[44] b[45] b[46] b[47] b[48]
+ b[49] b[4] b[50] b[51] b[52] b[53] b[54] b[55] b[56] b[57] b[58] b[59] b[5] b[60]
+ b[61] b[62] b[63] b[6] b[7] b[8] b[9] c[0] c[100] c[101] c[102] c[103] c[104] c[105]
+ c[106] c[107] c[108] c[109] c[10] c[110] c[111] c[112] c[113] c[114] c[115] c[116]
+ c[117] c[118] c[119] c[11] c[120] c[121] c[122] c[123] c[124] c[125] c[126] c[127]
+ c[12] c[13] c[14] c[15] c[16] c[17] c[18] c[19] c[1] c[20] c[21] c[22] c[23] c[24]
+ c[25] c[26] c[27] c[28] c[29] c[2] c[30] c[31] c[32] c[33] c[34] c[35] c[36] c[37]
+ c[38] c[39] c[3] c[40] c[41] c[42] c[43] c[44] c[45] c[46] c[47] c[48] c[49] c[4]
+ c[50] c[51] c[52] c[53] c[54] c[55] c[56] c[57] c[58] c[59] c[5] c[60] c[61] c[62]
+ c[63] c[64] c[65] c[66] c[67] c[68] c[69] c[6] c[70] c[71] c[72] c[73] c[74] c[75]
+ c[76] c[77] c[78] c[79] c[7] c[80] c[81] c[82] c[83] c[84] c[85] c[86] c[87] c[88]
+ c[89] c[8] c[90] c[91] c[92] c[93] c[94] c[95] c[96] c[97] c[98] c[99] c[9] clk
+ o[0] o[100] o[101] o[102] o[103] o[104] o[105] o[106] o[107] o[108] o[109] o[10]
+ o[110] o[111] o[112] o[113] o[114] o[115] o[116] o[117] o[118] o[119] o[11] o[120]
+ o[121] o[122] o[123] o[124] o[125] o[126] o[127] o[12] o[13] o[14] o[15] o[16] o[17]
+ o[18] o[19] o[1] o[20] o[21] o[22] o[23] o[24] o[25] o[26] o[27] o[28] o[29] o[2]
+ o[30] o[31] o[32] o[33] o[34] o[35] o[36] o[37] o[38] o[39] o[3] o[40] o[41] o[42]
+ o[43] o[44] o[45] o[46] o[47] o[48] o[49] o[4] o[50] o[51] o[52] o[53] o[54] o[55]
+ o[56] o[57] o[58] o[59] o[5] o[60] o[61] o[62] o[63] o[64] o[65] o[66] o[67] o[68]
+ o[69] o[6] o[70] o[71] o[72] o[73] o[74] o[75] o[76] o[77] o[78] o[79] o[7] o[80]
+ o[81] o[82] o[83] o[84] o[85] o[86] o[87] o[88] o[89] o[8] o[90] o[91] o[92] o[93]
+ o[94] o[95] o[96] o[97] o[98] o[99] o[9] rst
XFILLER_140_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_57_8 dadda_fa_1_57_8/A dadda_fa_1_57_8/B dadda_fa_1_57_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_58_3/A dadda_fa_3_57_0/A sky130_fd_sc_hd__fa_2
XFILLER_55_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_104_0 dadda_fa_2_104_0/A U$$2875/X U$$3008/X VGND VGND VPWR VPWR dadda_fa_3_105_2/CIN
+ dadda_fa_3_104_3/B sky130_fd_sc_hd__fa_1
XFILLER_63_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1290 U$$1290/A U$$1332/B VGND VGND VPWR VPWR U$$1290/X sky130_fd_sc_hd__xor2_1
XFILLER_10_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4244_1765 VGND VGND VPWR VPWR U$$4244_1765/HI U$$4244/B1 sky130_fd_sc_hd__conb_1
XFILLER_149_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_90_2 U$$2581/X U$$2714/X U$$2847/X VGND VGND VPWR VPWR dadda_fa_2_91_4/CIN
+ dadda_fa_2_90_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_85_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_282 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_83_1 U$$1769/X U$$1902/X U$$2035/X VGND VGND VPWR VPWR dadda_fa_2_84_2/A
+ dadda_fa_2_83_4/B sky130_fd_sc_hd__fa_1
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_60_0 dadda_fa_4_60_0/A dadda_fa_4_60_0/B dadda_fa_4_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/A dadda_fa_5_60_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_76_0 U$$1489/X U$$1622/X U$$1755/X VGND VGND VPWR VPWR dadda_fa_2_77_0/B
+ dadda_fa_2_76_3/B sky130_fd_sc_hd__fa_1
XFILLER_104_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3609 U$$3609/A U$$3609/B VGND VGND VPWR VPWR U$$3609/X sky130_fd_sc_hd__xor2_1
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2908 U$$2908/A U$$2988/B VGND VGND VPWR VPWR U$$2908/X sky130_fd_sc_hd__xor2_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_202 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_501_ _503_/CLK _501_/D VGND VGND VPWR VPWR _501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2919 U$$3193/A1 U$$2943/A2 U$$3056/B1 U$$2943/B2 VGND VGND VPWR VPWR U$$2920/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_213 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_5_124_1 U$$4511/X input156/X VGND VGND VPWR VPWR dadda_fa_6_125_0/CIN dadda_fa_7_124_0/A
+ sky130_fd_sc_hd__ha_1
XANTENNA_224 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _189_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 _194_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_432_ _432_/CLK _432_/D VGND VGND VPWR VPWR _432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_279 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_363_ _492_/CLK _363_/D VGND VGND VPWR VPWR _363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_294_ _615_/CLK _294_/D VGND VGND VPWR VPWR _294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_98_1 dadda_fa_3_98_1/A dadda_fa_3_98_1/B dadda_fa_3_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_0/CIN dadda_fa_4_98_2/A sky130_fd_sc_hd__fa_1
XFILLER_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_75_0 dadda_fa_6_75_0/A dadda_fa_6_75_0/B dadda_fa_6_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_76_0/B dadda_fa_7_75_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_5_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$370 U$$916/B1 U$$384/A2 U$$781/B1 U$$384/B2 VGND VGND VPWR VPWR U$$371/A sky130_fd_sc_hd__a22o_1
XU$$381 U$$381/A U$$383/B VGND VGND VPWR VPWR U$$381/X sky130_fd_sc_hd__xor2_1
XFILLER_178_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$392 U$$392/A1 U$$392/A2 U$$942/A1 U$$392/B2 VGND VGND VPWR VPWR U$$393/A sky130_fd_sc_hd__a22o_1
XFILLER_205_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_93_0 U$$2853/X U$$2986/X U$$3119/X VGND VGND VPWR VPWR dadda_fa_3_94_0/B
+ dadda_fa_3_93_2/B sky130_fd_sc_hd__fa_1
XFILLER_161_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1270 U$$3404/A1 VGND VGND VPWR VPWR U$$2171/A1 sky130_fd_sc_hd__buf_6
XFILLER_99_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1281 _605_/Q VGND VGND VPWR VPWR U$$3539/A1 sky130_fd_sc_hd__buf_4
Xrepeater1292 _603_/Q VGND VGND VPWR VPWR U$$3124/A1 sky130_fd_sc_hd__buf_4
XFILLER_141_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_62_6 dadda_fa_1_62_6/A dadda_fa_1_62_6/B dadda_fa_1_62_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_2/B dadda_fa_2_62_5/B sky130_fd_sc_hd__fa_1
XFILLER_45_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_55_5 U$$2777/X U$$2910/X U$$3043/X VGND VGND VPWR VPWR dadda_fa_2_56_2/A
+ dadda_fa_2_55_5/A sky130_fd_sc_hd__fa_1
XFILLER_110_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_48_4 U$$1699/X U$$1832/X U$$1965/X VGND VGND VPWR VPWR dadda_fa_2_49_2/B
+ dadda_fa_2_48_5/A sky130_fd_sc_hd__fa_1
XFILLER_167_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_18_2 dadda_fa_4_18_2/A dadda_fa_4_18_2/B dadda_ha_3_18_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_19_0/CIN dadda_fa_5_18_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_196_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_92_0 dadda_fa_7_92_0/A dadda_fa_7_92_0/B dadda_fa_7_92_0/CIN VGND VGND
+ VPWR VPWR _517_/D _388_/D sky130_fd_sc_hd__fa_2
XFILLER_17_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4107 U$$4516/B1 U$$4107/A2 U$$4107/B1 U$$4107/B2 VGND VGND VPWR VPWR U$$4108/A
+ sky130_fd_sc_hd__a22o_1
XU$$4118 U$$4392/A1 U$$4140/A2 U$$4394/A1 U$$4140/B2 VGND VGND VPWR VPWR U$$4119/A
+ sky130_fd_sc_hd__a22o_1
XU$$4129 U$$4129/A U$$4239/B VGND VGND VPWR VPWR U$$4129/X sky130_fd_sc_hd__xor2_1
XFILLER_59_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_670 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3406 U$$3952/B1 U$$3408/A2 U$$4504/A1 U$$3408/B2 VGND VGND VPWR VPWR U$$3407/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3417 U$$3417/A U$$3423/B VGND VGND VPWR VPWR U$$3417/X sky130_fd_sc_hd__xor2_1
XFILLER_19_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_394 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3428 _667_/Q U$$3428/B VGND VGND VPWR VPWR U$$3428/X sky130_fd_sc_hd__and2_1
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3439 U$$3713/A1 U$$3519/A2 U$$3578/A1 U$$3519/B2 VGND VGND VPWR VPWR U$$3440/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2705 U$$2705/A1 U$$2705/A2 U$$4214/A1 U$$2705/B2 VGND VGND VPWR VPWR U$$2706/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2716 U$$2716/A U$$2734/B VGND VGND VPWR VPWR U$$2716/X sky130_fd_sc_hd__xor2_1
XU$$2727 _610_/Q U$$2729/A2 _611_/Q U$$2729/B2 VGND VGND VPWR VPWR U$$2728/A sky130_fd_sc_hd__a22o_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2738 U$$2738/A U$$2739/A VGND VGND VPWR VPWR U$$2738/X sky130_fd_sc_hd__xor2_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2749 U$$2749/A U$$2795/B VGND VGND VPWR VPWR U$$2749/X sky130_fd_sc_hd__xor2_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_2 U$$845/X U$$978/X U$$1111/X VGND VGND VPWR VPWR dadda_fa_4_21_1/A
+ dadda_fa_4_20_2/B sky130_fd_sc_hd__fa_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_415_ _547_/CLK _415_/D VGND VGND VPWR VPWR _415_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1072 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_346_ _475_/CLK _346_/D VGND VGND VPWR VPWR _346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_277_ _523_/CLK _277_/D VGND VGND VPWR VPWR _277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_72_5 dadda_fa_2_72_5/A dadda_fa_2_72_5/B dadda_fa_2_72_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_2/A dadda_fa_4_72_0/A sky130_fd_sc_hd__fa_1
XFILLER_111_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_65_4 dadda_fa_2_65_4/A dadda_fa_2_65_4/B dadda_fa_2_65_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/CIN dadda_fa_3_65_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater904 _679_/Q VGND VGND VPWR VPWR U$$4296/B sky130_fd_sc_hd__buf_8
Xrepeater915 U$$4246/A VGND VGND VPWR VPWR U$$4239/B sky130_fd_sc_hd__buf_6
XFILLER_99_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater926 U$$4072/B VGND VGND VPWR VPWR U$$4084/B sky130_fd_sc_hd__clkbuf_8
XFILLER_83_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater937 U$$3943/B VGND VGND VPWR VPWR U$$3935/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_58_3 dadda_fa_2_58_3/A dadda_fa_2_58_3/B dadda_fa_2_58_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/B dadda_fa_3_58_3/B sky130_fd_sc_hd__fa_1
XFILLER_209_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater948 U$$3609/B VGND VGND VPWR VPWR U$$3613/B sky130_fd_sc_hd__buf_6
Xrepeater959 _667_/Q VGND VGND VPWR VPWR U$$3556/B sky130_fd_sc_hd__buf_6
Xdadda_fa_5_28_1 dadda_fa_5_28_1/A dadda_fa_5_28_1/B dadda_fa_5_28_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_29_0/B dadda_fa_7_28_0/A sky130_fd_sc_hd__fa_2
XU$$3940 U$$4214/A1 U$$3840/X U$$3942/A1 U$$3841/X VGND VGND VPWR VPWR U$$3941/A sky130_fd_sc_hd__a22o_1
XU$$3951 U$$3951/A U$$3973/A VGND VGND VPWR VPWR U$$3951/X sky130_fd_sc_hd__xor2_1
XU$$3962 U$$4236/A1 U$$3970/A2 U$$4238/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3963/A
+ sky130_fd_sc_hd__a22o_1
XU$$3973 U$$3973/A VGND VGND VPWR VPWR U$$3973/Y sky130_fd_sc_hd__inv_1
XU$$3984 U$$3984/A U$$3994/B VGND VGND VPWR VPWR U$$3984/X sky130_fd_sc_hd__xor2_1
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3995 U$$4269/A1 U$$4095/A2 _560_/Q U$$4105/B2 VGND VGND VPWR VPWR U$$3996/A sky130_fd_sc_hd__a22o_1
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_812 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_102_1 dadda_fa_5_102_1/A dadda_fa_5_102_1/B dadda_fa_5_102_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_103_0/B dadda_fa_7_102_0/A sky130_fd_sc_hd__fa_2
XFILLER_174_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput264 _274_/Q VGND VGND VPWR VPWR o[106] sky130_fd_sc_hd__buf_2
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput275 _284_/Q VGND VGND VPWR VPWR o[116] sky130_fd_sc_hd__buf_2
XFILLER_173_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3705_1755 VGND VGND VPWR VPWR U$$3705_1755/HI U$$3705/A1 sky130_fd_sc_hd__conb_1
XFILLER_160_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput286 _294_/Q VGND VGND VPWR VPWR o[126] sky130_fd_sc_hd__buf_2
XFILLER_87_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput297 _188_/Q VGND VGND VPWR VPWR o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_60_3 U$$3186/X U$$3319/X U$$3452/X VGND VGND VPWR VPWR dadda_fa_2_61_1/B
+ dadda_fa_2_60_4/B sky130_fd_sc_hd__fa_1
XFILLER_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_2 U$$1177/X U$$1310/X U$$1443/X VGND VGND VPWR VPWR dadda_fa_2_54_1/A
+ dadda_fa_2_53_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_30_1 dadda_fa_4_30_1/A dadda_fa_4_30_1/B dadda_fa_4_30_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/B dadda_fa_5_30_1/B sky130_fd_sc_hd__fa_1
XFILLER_28_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_46_1 U$$498/X U$$631/X U$$764/X VGND VGND VPWR VPWR dadda_fa_2_47_2/A
+ dadda_fa_2_46_4/B sky130_fd_sc_hd__fa_1
XFILLER_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_23_0 dadda_fa_4_23_0/A dadda_fa_4_23_0/B dadda_fa_4_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/A dadda_fa_5_23_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_39_0 U$$85/X U$$218/X U$$351/X VGND VGND VPWR VPWR dadda_fa_2_40_4/A dadda_fa_2_39_5/B
+ sky130_fd_sc_hd__fa_1
XFILLER_208_1020 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_200_ _478_/CLK _200_/D VGND VGND VPWR VPWR _200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_75_3 dadda_fa_3_75_3/A dadda_fa_3_75_3/B dadda_fa_3_75_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_1/B dadda_fa_4_75_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_68_2 dadda_fa_3_68_2/A dadda_fa_3_68_2/B dadda_fa_3_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_1/A dadda_fa_4_68_2/B sky130_fd_sc_hd__fa_1
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_38_0 dadda_fa_6_38_0/A dadda_fa_6_38_0/B dadda_fa_6_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_39_0/B dadda_fa_7_38_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3203 _574_/Q U$$3285/A2 _575_/Q U$$3285/B2 VGND VGND VPWR VPWR U$$3204/A sky130_fd_sc_hd__a22o_1
XU$$3214 U$$3214/A U$$3218/B VGND VGND VPWR VPWR U$$3214/X sky130_fd_sc_hd__xor2_1
XFILLER_24_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3225 U$$4184/A1 U$$3273/A2 U$$4186/A1 U$$3273/B2 VGND VGND VPWR VPWR U$$3226/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3236 U$$3236/A U$$3236/B VGND VGND VPWR VPWR U$$3236/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2502 U$$2774/B1 U$$2550/A2 U$$2641/A1 U$$2550/B2 VGND VGND VPWR VPWR U$$2503/A
+ sky130_fd_sc_hd__a22o_1
XU$$3247 U$$3932/A1 U$$3273/A2 U$$918/B1 U$$3273/B2 VGND VGND VPWR VPWR U$$3248/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$18 _442_/Q _314_/Q VGND VGND VPWR VPWR final_adder.U$$513/B1 final_adder.U$$640/A
+ sky130_fd_sc_hd__ha_2
XU$$3258 U$$3258/A U$$3272/B VGND VGND VPWR VPWR U$$3258/X sky130_fd_sc_hd__xor2_1
XU$$2513 U$$2513/A U$$2551/B VGND VGND VPWR VPWR U$$2513/X sky130_fd_sc_hd__xor2_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$29 _453_/Q _325_/Q VGND VGND VPWR VPWR final_adder.U$$157/B1 final_adder.U$$651/A
+ sky130_fd_sc_hd__ha_2
XFILLER_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2524 U$$2796/B1 U$$2524/A2 U$$334/A1 U$$2524/B2 VGND VGND VPWR VPWR U$$2525/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3269 U$$3952/B1 U$$3273/A2 U$$3269/B1 U$$3273/B2 VGND VGND VPWR VPWR U$$3270/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2535 U$$2535/A _653_/Q VGND VGND VPWR VPWR U$$2535/X sky130_fd_sc_hd__xor2_1
XU$$1801 U$$2210/B1 U$$1851/A2 U$$20/B1 U$$1851/B2 VGND VGND VPWR VPWR U$$1802/A sky130_fd_sc_hd__a22o_1
XU$$2546 U$$900/B1 U$$2566/A2 U$$3096/A1 U$$2566/B2 VGND VGND VPWR VPWR U$$2547/A
+ sky130_fd_sc_hd__a22o_1
XU$$2557 U$$2557/A U$$2597/B VGND VGND VPWR VPWR U$$2557/X sky130_fd_sc_hd__xor2_1
XU$$1812 U$$1812/A U$$1852/B VGND VGND VPWR VPWR U$$1812/X sky130_fd_sc_hd__xor2_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2568 U$$4075/A1 U$$2580/A2 U$$4351/A1 U$$2580/B2 VGND VGND VPWR VPWR U$$2569/A
+ sky130_fd_sc_hd__a22o_1
XU$$1823 U$$999/B1 U$$1855/A2 U$$866/A1 U$$1855/B2 VGND VGND VPWR VPWR U$$1824/A sky130_fd_sc_hd__a22o_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1834 U$$1834/A U$$1852/B VGND VGND VPWR VPWR U$$1834/X sky130_fd_sc_hd__xor2_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2579 U$$2579/A U$$2583/B VGND VGND VPWR VPWR U$$2579/X sky130_fd_sc_hd__xor2_1
XU$$1845 U$$3352/A1 U$$1897/A2 U$$3217/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1846/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1856 U$$1856/A U$$1874/B VGND VGND VPWR VPWR U$$1856/X sky130_fd_sc_hd__xor2_1
XU$$1867 U$$3374/A1 U$$1785/X U$$2963/B1 U$$1786/X VGND VGND VPWR VPWR U$$1868/A sky130_fd_sc_hd__a22o_1
XFILLER_199_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1878 U$$1878/A U$$1884/B VGND VGND VPWR VPWR U$$1878/X sky130_fd_sc_hd__xor2_1
XU$$1889 U$$3122/A1 U$$1897/A2 U$$3124/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1890/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_329_ _458_/CLK _329_/D VGND VGND VPWR VPWR _329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_70_2 dadda_fa_2_70_2/A dadda_fa_2_70_2/B dadda_fa_2_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/A dadda_fa_3_70_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_63_1 dadda_fa_2_63_1/A dadda_fa_2_63_1/B dadda_fa_2_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_0/CIN dadda_fa_3_63_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater701 U$$4071/B2 VGND VGND VPWR VPWR U$$4061/B2 sky130_fd_sc_hd__buf_4
XFILLER_96_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater712 U$$3823/B2 VGND VGND VPWR VPWR U$$3833/B2 sky130_fd_sc_hd__buf_4
Xrepeater723 U$$3664/B2 VGND VGND VPWR VPWR U$$3662/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_5_40_0 dadda_fa_5_40_0/A dadda_fa_5_40_0/B dadda_fa_5_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_41_0/A dadda_fa_6_40_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$519 final_adder.U$$646/A final_adder.U$$646/B final_adder.U$$519/B1
+ VGND VGND VPWR VPWR final_adder.U$$647/B sky130_fd_sc_hd__a21o_1
Xdadda_fa_2_56_0 dadda_fa_2_56_0/A dadda_fa_2_56_0/B dadda_fa_2_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_0/B dadda_fa_3_56_2/B sky130_fd_sc_hd__fa_1
Xrepeater734 U$$3418/B2 VGND VGND VPWR VPWR U$$3368/B2 sky130_fd_sc_hd__buf_6
Xrepeater745 U$$3283/B2 VGND VGND VPWR VPWR U$$3231/B2 sky130_fd_sc_hd__buf_6
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater756 U$$3144/B2 VGND VGND VPWR VPWR U$$3132/B2 sky130_fd_sc_hd__buf_4
XFILLER_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater767 U$$308/B2 VGND VGND VPWR VPWR U$$318/B2 sky130_fd_sc_hd__buf_4
Xrepeater778 U$$2745/X VGND VGND VPWR VPWR U$$2798/B2 sky130_fd_sc_hd__buf_4
XU$$4460 _586_/Q U$$4388/X _587_/Q U$$4468/B2 VGND VGND VPWR VPWR U$$4461/A sky130_fd_sc_hd__a22o_1
XFILLER_38_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4471 U$$4471/A U$$4471/B VGND VGND VPWR VPWR U$$4471/X sky130_fd_sc_hd__xor2_1
Xrepeater789 U$$2608/X VGND VGND VPWR VPWR U$$2733/B2 sky130_fd_sc_hd__buf_4
XU$$4482 U$$4482/A1 U$$4388/X U$$4484/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4483/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4493 U$$4493/A U$$4493/B VGND VGND VPWR VPWR U$$4493/X sky130_fd_sc_hd__xor2_1
XU$$3770 U$$3770/A U$$3816/B VGND VGND VPWR VPWR U$$3770/X sky130_fd_sc_hd__xor2_1
XU$$3781 U$$4466/A1 U$$3795/A2 U$$4468/A1 U$$3795/B2 VGND VGND VPWR VPWR U$$3782/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3792 U$$3792/A U$$3804/B VGND VGND VPWR VPWR U$$3792/X sky130_fd_sc_hd__xor2_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1040 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_85_2 dadda_fa_4_85_2/A dadda_fa_4_85_2/B dadda_fa_4_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/CIN dadda_fa_5_85_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_78_1 dadda_fa_4_78_1/A dadda_fa_4_78_1/B dadda_fa_4_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/B dadda_fa_5_78_1/B sky130_fd_sc_hd__fa_1
XFILLER_134_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_55_0 dadda_fa_7_55_0/A dadda_fa_7_55_0/B dadda_fa_7_55_0/CIN VGND VGND
+ VPWR VPWR _480_/D _351_/D sky130_fd_sc_hd__fa_1
XFILLER_134_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$903 U$$903/A U$$907/B VGND VGND VPWR VPWR U$$903/X sky130_fd_sc_hd__xor2_1
XFILLER_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$914 U$$914/A1 U$$956/A2 U$$914/B1 U$$956/B2 VGND VGND VPWR VPWR U$$915/A sky130_fd_sc_hd__a22o_1
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$925 U$$925/A U$$925/B VGND VGND VPWR VPWR U$$925/X sky130_fd_sc_hd__xor2_1
XU$$936 U$$936/A1 U$$826/X U$$938/A1 U$$827/X VGND VGND VPWR VPWR U$$937/A sky130_fd_sc_hd__a22o_1
XFILLER_84_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$947 U$$947/A U$$951/B VGND VGND VPWR VPWR U$$947/X sky130_fd_sc_hd__xor2_1
XU$$958 U$$958/A VGND VGND VPWR VPWR U$$958/Y sky130_fd_sc_hd__inv_1
XU$$969 U$$969/A1 U$$995/A2 U$$971/A1 U$$995/B2 VGND VGND VPWR VPWR U$$970/A sky130_fd_sc_hd__a22o_1
XU$$1108 U$$695/B1 U$$1150/A2 U$$562/A1 U$$1150/B2 VGND VGND VPWR VPWR U$$1109/A sky130_fd_sc_hd__a22o_1
XU$$1119 U$$1119/A U$$1151/B VGND VGND VPWR VPWR U$$1119/X sky130_fd_sc_hd__xor2_1
XFILLER_71_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1072 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1064 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_80_1 dadda_fa_3_80_1/A dadda_fa_3_80_1/B dadda_fa_3_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_0/CIN dadda_fa_4_80_2/A sky130_fd_sc_hd__fa_1
XFILLER_152_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_73_0 dadda_fa_3_73_0/A dadda_fa_3_73_0/B dadda_fa_3_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_0/B dadda_fa_4_73_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3000 U$$3000/A U$$3000/B VGND VGND VPWR VPWR U$$3000/X sky130_fd_sc_hd__xor2_1
XU$$3011 U$$3285/A1 U$$2881/X U$$3011/B1 U$$2882/X VGND VGND VPWR VPWR U$$3012/A sky130_fd_sc_hd__a22o_1
XU$$3022 U$$3157/B1 U$$3054/A2 U$$3022/B1 U$$3054/B2 VGND VGND VPWR VPWR U$$3023/A
+ sky130_fd_sc_hd__a22o_1
XU$$3033 U$$3033/A U$$3049/B VGND VGND VPWR VPWR U$$3033/X sky130_fd_sc_hd__xor2_1
XFILLER_75_971 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3044 U$$4140/A1 U$$3082/A2 U$$3181/B1 U$$3082/B2 VGND VGND VPWR VPWR U$$3045/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3055 U$$3055/A U$$3065/B VGND VGND VPWR VPWR U$$3055/X sky130_fd_sc_hd__xor2_1
XU$$2310 U$$4502/A1 U$$2318/A2 U$$940/B1 U$$2318/B2 VGND VGND VPWR VPWR U$$2311/A
+ sky130_fd_sc_hd__a22o_1
XU$$2321 U$$2321/A U$$2321/B VGND VGND VPWR VPWR U$$2321/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_5 U$$2338/X input185/X dadda_fa_2_35_5/CIN VGND VGND VPWR VPWR dadda_fa_3_36_2/A
+ dadda_fa_4_35_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_102_0 dadda_fa_4_102_0/A dadda_fa_4_102_0/B dadda_fa_4_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/A dadda_fa_5_102_1/A sky130_fd_sc_hd__fa_1
XU$$3066 U$$4436/A1 U$$3066/A2 U$$4436/B1 U$$3066/B2 VGND VGND VPWR VPWR U$$3067/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2332 U$$2466/A U$$2332/B VGND VGND VPWR VPWR U$$2332/X sky130_fd_sc_hd__and2_1
XU$$3077 U$$3077/A U$$3077/B VGND VGND VPWR VPWR U$$3077/X sky130_fd_sc_hd__xor2_1
XU$$2343 U$$2343/A1 U$$2367/A2 U$$2345/A1 U$$2367/B2 VGND VGND VPWR VPWR U$$2344/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3088 U$$3088/A1 U$$3120/A2 U$$4186/A1 U$$3120/B2 VGND VGND VPWR VPWR U$$3089/A
+ sky130_fd_sc_hd__a22o_1
XU$$2354 U$$2354/A U$$2400/B VGND VGND VPWR VPWR U$$2354/X sky130_fd_sc_hd__xor2_1
XU$$3099 U$$3099/A U$$3111/B VGND VGND VPWR VPWR U$$3099/X sky130_fd_sc_hd__xor2_1
XU$$1620 U$$1620/A U$$1628/B VGND VGND VPWR VPWR U$$1620/X sky130_fd_sc_hd__xor2_1
XU$$2365 U$$582/B1 U$$2367/A2 U$$449/A1 U$$2367/B2 VGND VGND VPWR VPWR U$$2366/A sky130_fd_sc_hd__a22o_1
XFILLER_201_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2376 U$$2376/A U$$2418/B VGND VGND VPWR VPWR U$$2376/X sky130_fd_sc_hd__xor2_1
XU$$1631 U$$2314/B1 U$$1635/A2 U$$2866/A1 U$$1635/B2 VGND VGND VPWR VPWR U$$1632/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1642 U$$1642/A U$$1642/B VGND VGND VPWR VPWR U$$1642/X sky130_fd_sc_hd__xor2_1
XFILLER_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2387 U$$467/B1 U$$2387/A2 U$$334/A1 U$$2387/B2 VGND VGND VPWR VPWR U$$2388/A sky130_fd_sc_hd__a22o_1
XFILLER_76_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2398 U$$2398/A U$$2442/B VGND VGND VPWR VPWR U$$2398/X sky130_fd_sc_hd__xor2_1
XU$$1653 U$$1653/A U$$1687/B VGND VGND VPWR VPWR U$$1653/X sky130_fd_sc_hd__xor2_1
XU$$4381_1767 VGND VGND VPWR VPWR U$$4381_1767/HI U$$4381/B1 sky130_fd_sc_hd__conb_1
XU$$1664 U$$840/B1 U$$1684/A2 U$$568/B1 U$$1684/B2 VGND VGND VPWR VPWR U$$1665/A sky130_fd_sc_hd__a22o_1
XFILLER_163_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1675 U$$1675/A U$$1711/B VGND VGND VPWR VPWR U$$1675/X sky130_fd_sc_hd__xor2_1
XU$$1686 U$$42/A1 U$$1736/A2 U$$42/B1 U$$1736/B2 VGND VGND VPWR VPWR U$$1687/A sky130_fd_sc_hd__a22o_1
XFILLER_163_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1697 U$$1697/A U$$1723/B VGND VGND VPWR VPWR U$$1697/X sky130_fd_sc_hd__xor2_1
XFILLER_202_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_95_1 dadda_fa_5_95_1/A dadda_fa_5_95_1/B dadda_fa_5_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_96_0/B dadda_fa_7_95_0/A sky130_fd_sc_hd__fa_1
XFILLER_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_88_0 dadda_fa_5_88_0/A dadda_fa_5_88_0/B dadda_fa_5_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_89_0/A dadda_fa_6_88_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_200_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$305 final_adder.U$$304/A final_adder.U$$225/X final_adder.U$$227/X
+ VGND VGND VPWR VPWR final_adder.U$$305/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$316 final_adder.U$$316/A final_adder.U$$316/B VGND VGND VPWR VPWR
+ final_adder.U$$316/X sky130_fd_sc_hd__and2_1
Xrepeater520 U$$334/A2 VGND VGND VPWR VPWR U$$308/A2 sky130_fd_sc_hd__buf_4
Xrepeater531 U$$2744/X VGND VGND VPWR VPWR U$$2832/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$327 final_adder.U$$326/A final_adder.U$$269/X final_adder.U$$271/X
+ VGND VGND VPWR VPWR final_adder.U$$327/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$338 final_adder.U$$338/A final_adder.U$$338/B VGND VGND VPWR VPWR
+ final_adder.U$$360/A sky130_fd_sc_hd__and2_1
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater542 U$$2607/X VGND VGND VPWR VPWR U$$2707/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$349 final_adder.U$$348/A final_adder.U$$313/X final_adder.U$$315/X
+ VGND VGND VPWR VPWR final_adder.U$$349/X sky130_fd_sc_hd__a21o_1
XFILLER_38_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater553 U$$2395/A2 VGND VGND VPWR VPWR U$$2387/A2 sky130_fd_sc_hd__buf_6
Xrepeater564 U$$2196/X VGND VGND VPWR VPWR U$$2274/A2 sky130_fd_sc_hd__buf_4
Xrepeater575 U$$2040/A2 VGND VGND VPWR VPWR U$$1956/A2 sky130_fd_sc_hd__buf_6
Xrepeater586 U$$1907/A2 VGND VGND VPWR VPWR U$$1855/A2 sky130_fd_sc_hd__buf_8
XFILLER_77_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater597 U$$1778/A2 VGND VGND VPWR VPWR U$$1740/A2 sky130_fd_sc_hd__buf_12
XFILLER_84_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4290 U$$4290/A U$$4296/B VGND VGND VPWR VPWR U$$4290/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_90_0 dadda_fa_4_90_0/A dadda_fa_4_90_0/B dadda_fa_4_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/A dadda_fa_5_90_1/A sky130_fd_sc_hd__fa_1
XFILLER_107_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1043 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_104_2 input134/X dadda_fa_3_104_2/B dadda_fa_3_104_2/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_105_1/A dadda_fa_4_104_2/B sky130_fd_sc_hd__fa_1
XFILLER_122_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_118_0 dadda_fa_6_118_0/A dadda_fa_6_118_0/B dadda_fa_6_118_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_119_0/B dadda_fa_7_118_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$700 U$$700/A U$$726/B VGND VGND VPWR VPWR U$$700/X sky130_fd_sc_hd__xor2_1
X_663_ _674_/CLK _663_/D VGND VGND VPWR VPWR _663_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$711 U$$848/A1 U$$765/A2 U$$848/B1 U$$765/B2 VGND VGND VPWR VPWR U$$712/A sky130_fd_sc_hd__a22o_1
XFILLER_90_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_38_3 dadda_fa_3_38_3/A dadda_fa_3_38_3/B dadda_fa_3_38_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_1/B dadda_fa_4_38_2/CIN sky130_fd_sc_hd__fa_1
XU$$722 U$$722/A U$$760/B VGND VGND VPWR VPWR U$$722/X sky130_fd_sc_hd__xor2_1
XFILLER_75_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$733 U$$733/A1 U$$759/A2 U$$733/B1 U$$759/B2 VGND VGND VPWR VPWR U$$734/A sky130_fd_sc_hd__a22o_1
XFILLER_205_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$744 U$$744/A U$$748/B VGND VGND VPWR VPWR U$$744/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_594_ _596_/CLK _594_/D VGND VGND VPWR VPWR _594_/Q sky130_fd_sc_hd__dfxtp_2
XU$$755 U$$890/B1 U$$795/A2 U$$757/A1 U$$795/B2 VGND VGND VPWR VPWR U$$756/A sky130_fd_sc_hd__a22o_1
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$766 U$$766/A U$$766/B VGND VGND VPWR VPWR U$$766/X sky130_fd_sc_hd__xor2_1
XU$$777 U$$912/B1 U$$783/A2 U$$914/B1 U$$783/B2 VGND VGND VPWR VPWR U$$778/A sky130_fd_sc_hd__a22o_1
XU$$788 U$$788/A U$$810/B VGND VGND VPWR VPWR U$$788/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$799 U$$936/A1 U$$689/X U$$938/A1 U$$690/X VGND VGND VPWR VPWR U$$800/A sky130_fd_sc_hd__a22o_1
XFILLER_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1600 U$$4418/A1 VGND VGND VPWR VPWR U$$2909/B1 sky130_fd_sc_hd__buf_6
XFILLER_126_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1611 _564_/Q VGND VGND VPWR VPWR U$$4416/A1 sky130_fd_sc_hd__buf_6
XANTENNA_5 _456_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1622 U$$987/A1 VGND VGND VPWR VPWR U$$302/A1 sky130_fd_sc_hd__buf_6
XFILLER_67_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1633 U$$4273/A1 VGND VGND VPWR VPWR U$$4136/A1 sky130_fd_sc_hd__buf_6
Xrepeater1644 U$$3447/B1 VGND VGND VPWR VPWR U$$4408/A1 sky130_fd_sc_hd__buf_6
XFILLER_67_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1655 U$$429/B1 VGND VGND VPWR VPWR U$$20/A1 sky130_fd_sc_hd__buf_6
Xrepeater1666 U$$2893/B1 VGND VGND VPWR VPWR U$$429/A1 sky130_fd_sc_hd__buf_4
XFILLER_98_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1677 U$$3713/B1 VGND VGND VPWR VPWR U$$3578/A1 sky130_fd_sc_hd__buf_6
XFILLER_113_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1688 U$$2613/B1 VGND VGND VPWR VPWR U$$695/B1 sky130_fd_sc_hd__buf_4
XFILLER_99_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1699 U$$556/B1 VGND VGND VPWR VPWR U$$2611/B1 sky130_fd_sc_hd__buf_6
XFILLER_112_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_40_3 U$$2747/X U$$2787/B input191/X VGND VGND VPWR VPWR dadda_fa_3_41_1/B
+ dadda_fa_3_40_3/B sky130_fd_sc_hd__fa_1
XFILLER_94_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_33_2 U$$871/X U$$1004/X U$$1137/X VGND VGND VPWR VPWR dadda_fa_3_34_1/A
+ dadda_fa_3_33_3/A sky130_fd_sc_hd__fa_1
XFILLER_207_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2140 U$$2140/A U$$2174/B VGND VGND VPWR VPWR U$$2140/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_10_1 dadda_fa_5_10_1/A dadda_fa_5_10_1/B dadda_ha_4_10_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_11_0/B dadda_fa_7_10_0/A sky130_fd_sc_hd__fa_1
XU$$2151 U$$3519/B1 U$$2189/A2 U$$781/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2152/A
+ sky130_fd_sc_hd__a22o_1
XU$$2162 U$$2162/A U$$2170/B VGND VGND VPWR VPWR U$$2162/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_26_1 U$$458/X U$$591/X U$$724/X VGND VGND VPWR VPWR dadda_fa_3_27_2/CIN
+ dadda_fa_3_26_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2173 U$$940/A1 U$$2059/X U$$4228/B1 U$$2060/X VGND VGND VPWR VPWR U$$2174/A sky130_fd_sc_hd__a22o_1
XU$$2184 U$$2184/A U$$2186/B VGND VGND VPWR VPWR U$$2184/X sky130_fd_sc_hd__xor2_1
XFILLER_23_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1450 U$$900/B1 U$$1478/A2 U$$3096/A1 U$$1478/B2 VGND VGND VPWR VPWR U$$1451/A
+ sky130_fd_sc_hd__a22o_1
XU$$2195 _649_/Q U$$2195/B VGND VGND VPWR VPWR U$$2195/X sky130_fd_sc_hd__and2_1
XU$$1461 U$$1461/A U$$1475/B VGND VGND VPWR VPWR U$$1461/X sky130_fd_sc_hd__xor2_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1472 U$$924/A1 U$$1474/A2 U$$924/B1 U$$1474/B2 VGND VGND VPWR VPWR U$$1473/A sky130_fd_sc_hd__a22o_1
XFILLER_50_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1483 U$$1483/A U$$1501/B VGND VGND VPWR VPWR U$$1483/X sky130_fd_sc_hd__xor2_1
XFILLER_194_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1494 U$$2588/B1 U$$1500/A2 U$$948/A1 U$$1500/B2 VGND VGND VPWR VPWR U$$1495/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_85_5 U$$3502/X U$$3635/X U$$3768/X VGND VGND VPWR VPWR dadda_fa_2_86_4/A
+ dadda_fa_3_85_0/A sky130_fd_sc_hd__fa_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_78_4 U$$2823/X U$$2956/X U$$3089/X VGND VGND VPWR VPWR dadda_fa_2_79_1/CIN
+ dadda_fa_2_78_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$102 _526_/Q _398_/Q VGND VGND VPWR VPWR final_adder.U$$597/B1 final_adder.U$$724/A
+ sky130_fd_sc_hd__ha_1
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$113 _537_/Q _409_/Q VGND VGND VPWR VPWR final_adder.U$$241/B1 final_adder.U$$735/A
+ sky130_fd_sc_hd__ha_2
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$124 _548_/Q _420_/Q VGND VGND VPWR VPWR final_adder.U$$619/B1 final_adder.U$$746/A
+ sky130_fd_sc_hd__ha_2
Xdadda_fa_4_48_2 dadda_fa_4_48_2/A dadda_fa_4_48_2/B dadda_fa_4_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/CIN dadda_fa_5_48_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$135 final_adder.U$$7/SUM final_adder.U$$6/COUT final_adder.U$$7/COUT
+ VGND VGND VPWR VPWR final_adder.U$$135/X sky130_fd_sc_hd__a21o_1
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$146 final_adder.U$$641/A final_adder.U$$640/A VGND VGND VPWR VPWR
+ final_adder.U$$264/A sky130_fd_sc_hd__and2_1
XFILLER_100_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_971 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$157 final_adder.U$$651/A final_adder.U$$523/B1 final_adder.U$$157/B1
+ VGND VGND VPWR VPWR final_adder.U$$157/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$168 final_adder.U$$663/A final_adder.U$$662/A VGND VGND VPWR VPWR
+ final_adder.U$$276/B sky130_fd_sc_hd__and2_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$179 final_adder.U$$673/A final_adder.U$$545/B1 final_adder.U$$179/B1
+ VGND VGND VPWR VPWR final_adder.U$$179/X sky130_fd_sc_hd__a21o_1
XFILLER_174_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater394 U$$826/X VGND VGND VPWR VPWR U$$928/A2 sky130_fd_sc_hd__buf_4
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_18_0 dadda_fa_7_18_0/A dadda_fa_7_18_0/B dadda_fa_7_18_0/CIN VGND VGND
+ VPWR VPWR _443_/D _314_/D sky130_fd_sc_hd__fa_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4405_1781 VGND VGND VPWR VPWR U$$4405_1781/HI U$$4405/B sky130_fd_sc_hd__conb_1
XFILLER_166_331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput120 b[5] VGND VGND VPWR VPWR _557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_209_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput131 c[101] VGND VGND VPWR VPWR input131/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_50_2 dadda_fa_3_50_2/A dadda_fa_3_50_2/B dadda_fa_3_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_1/A dadda_fa_4_50_2/B sky130_fd_sc_hd__fa_1
XFILLER_23_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput142 c[111] VGND VGND VPWR VPWR input142/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_1139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_66_2 U$$937/X U$$1070/X U$$1203/X VGND VGND VPWR VPWR dadda_fa_1_67_6/A
+ dadda_fa_1_66_8/A sky130_fd_sc_hd__fa_1
Xinput153 c[121] VGND VGND VPWR VPWR input153/X sky130_fd_sc_hd__clkbuf_1
XTAP_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput164 c[16] VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__clkbuf_1
XTAP_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 c[26] VGND VGND VPWR VPWR input175/X sky130_fd_sc_hd__clkbuf_2
XTAP_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 c[36] VGND VGND VPWR VPWR input186/X sky130_fd_sc_hd__buf_4
Xdadda_fa_3_43_1 dadda_fa_3_43_1/A dadda_fa_3_43_1/B dadda_fa_3_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_0/CIN dadda_fa_4_43_2/A sky130_fd_sc_hd__fa_1
XFILLER_91_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_59_1 U$$524/X U$$657/X U$$790/X VGND VGND VPWR VPWR dadda_fa_1_60_6/CIN
+ dadda_fa_1_59_8/B sky130_fd_sc_hd__fa_1
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput197 c[46] VGND VGND VPWR VPWR input197/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_20_0 dadda_fa_6_20_0/A dadda_fa_6_20_0/B dadda_fa_6_20_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_21_0/B dadda_fa_7_20_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$680 final_adder.U$$680/A final_adder.U$$680/B VGND VGND VPWR VPWR
+ _226_/D sky130_fd_sc_hd__xor2_1
XTAP_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_36_0 dadda_fa_3_36_0/A dadda_fa_3_36_0/B dadda_fa_3_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_0/B dadda_fa_4_36_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$530 U$$530/A U$$532/B VGND VGND VPWR VPWR U$$530/X sky130_fd_sc_hd__xor2_1
X_646_ _648_/CLK _646_/D VGND VGND VPWR VPWR _646_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$691 final_adder.U$$691/A final_adder.U$$691/B VGND VGND VPWR VPWR
+ _237_/D sky130_fd_sc_hd__xor2_4
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$541 U$$676/B1 U$$545/A2 U$$678/B1 U$$545/B2 VGND VGND VPWR VPWR U$$542/A sky130_fd_sc_hd__a22o_1
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$552 U$$550/Y _624_/Q _623_/Q U$$551/X U$$548/Y VGND VGND VPWR VPWR U$$552/X sky130_fd_sc_hd__a32o_2
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$563 U$$563/A U$$589/B VGND VGND VPWR VPWR U$$563/X sky130_fd_sc_hd__xor2_1
XU$$574 U$$26/A1 U$$574/A2 U$$28/A1 U$$574/B2 VGND VGND VPWR VPWR U$$575/A sky130_fd_sc_hd__a22o_1
X_577_ _582_/CLK _577_/D VGND VGND VPWR VPWR _577_/Q sky130_fd_sc_hd__dfxtp_4
XU$$585 U$$585/A U$$627/B VGND VGND VPWR VPWR U$$585/X sky130_fd_sc_hd__xor2_1
XU$$596 U$$596/A1 U$$622/A2 U$$596/B1 U$$622/B2 VGND VGND VPWR VPWR U$$597/A sky130_fd_sc_hd__a22o_1
XFILLER_71_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_95_4 U$$4187/X U$$4320/X U$$4453/X VGND VGND VPWR VPWR dadda_fa_3_96_1/CIN
+ dadda_fa_3_95_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1430 U$$4186/A1 VGND VGND VPWR VPWR U$$3362/B1 sky130_fd_sc_hd__buf_6
XFILLER_132_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1441 U$$4456/B1 VGND VGND VPWR VPWR U$$3771/B1 sky130_fd_sc_hd__buf_6
XFILLER_172_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3842_1757 VGND VGND VPWR VPWR U$$3842_1757/HI U$$3842/A1 sky130_fd_sc_hd__conb_1
Xrepeater1452 U$$3358/A1 VGND VGND VPWR VPWR U$$70/A1 sky130_fd_sc_hd__buf_4
Xrepeater1463 U$$4450/B1 VGND VGND VPWR VPWR U$$3354/B1 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_2_88_3 dadda_fa_2_88_3/A dadda_fa_2_88_3/B dadda_fa_2_88_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_1/B dadda_fa_3_88_3/B sky130_fd_sc_hd__fa_1
XFILLER_125_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1474 _581_/Q VGND VGND VPWR VPWR U$$4450/A1 sky130_fd_sc_hd__buf_6
Xrepeater1485 U$$334/B1 VGND VGND VPWR VPWR U$$62/A1 sky130_fd_sc_hd__buf_4
XFILLER_67_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1496 U$$4031/B1 VGND VGND VPWR VPWR U$$334/A1 sky130_fd_sc_hd__buf_6
XFILLER_99_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_58_1 dadda_fa_5_58_1/A dadda_fa_5_58_1/B dadda_fa_5_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_59_0/B dadda_fa_7_58_0/A sky130_fd_sc_hd__fa_2
XFILLER_80_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_104_1 U$$3141/X U$$3274/X U$$3407/X VGND VGND VPWR VPWR dadda_fa_3_105_3/A
+ dadda_fa_3_104_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1280 U$$1280/A U$$1280/B VGND VGND VPWR VPWR U$$1280/X sky130_fd_sc_hd__xor2_1
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1291 U$$467/B1 U$$1291/A2 U$$334/A1 U$$1291/B2 VGND VGND VPWR VPWR U$$1292/A sky130_fd_sc_hd__a22o_1
XFILLER_210_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_125_0 U$$4246/Y U$$4380/X U$$4513/X VGND VGND VPWR VPWR dadda_fa_6_126_0/CIN
+ dadda_fa_7_125_0/A sky130_fd_sc_hd__fa_1
XFILLER_149_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_83_2 U$$2168/X U$$2301/X U$$2434/X VGND VGND VPWR VPWR dadda_fa_2_84_2/B
+ dadda_fa_2_83_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_116_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_60_1 dadda_fa_4_60_1/A dadda_fa_4_60_1/B dadda_fa_4_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/B dadda_fa_5_60_1/B sky130_fd_sc_hd__fa_1
XFILLER_120_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_76_1 U$$1888/X U$$2021/X U$$2154/X VGND VGND VPWR VPWR dadda_fa_2_77_0/CIN
+ dadda_fa_2_76_3/CIN sky130_fd_sc_hd__fa_1
XU$$4435_1796 VGND VGND VPWR VPWR U$$4435_1796/HI U$$4435/B sky130_fd_sc_hd__conb_1
XFILLER_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_53_0 dadda_fa_4_53_0/A dadda_fa_4_53_0/B dadda_fa_4_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/A dadda_fa_5_53_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_69_0 U$$2406/X U$$2539/X U$$2672/X VGND VGND VPWR VPWR dadda_fa_2_70_0/B
+ dadda_fa_2_69_3/B sky130_fd_sc_hd__fa_1
XFILLER_86_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2909 U$$2909/A1 U$$2959/A2 U$$2909/B1 U$$2959/B2 VGND VGND VPWR VPWR U$$2910/A
+ sky130_fd_sc_hd__a22o_1
X_500_ _500_/CLK _500_/D VGND VGND VPWR VPWR _500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_214 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_225 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 _189_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_431_ _431_/CLK _431_/D VGND VGND VPWR VPWR _431_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_6__f_clk clkbuf_2_3_0_clk/X VGND VGND VPWR VPWR _369_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 _194_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_258 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_269 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_362_ _491_/CLK _362_/D VGND VGND VPWR VPWR _362_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_293_ _615_/CLK _293_/D VGND VGND VPWR VPWR _293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_114_0_1869 VGND VGND VPWR VPWR dadda_fa_3_114_0/A dadda_fa_3_114_0_1869/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_158_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_98_2 dadda_fa_3_98_2/A dadda_fa_3_98_2/B dadda_fa_3_98_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_1/A dadda_fa_4_98_2/B sky130_fd_sc_hd__fa_1
XFILLER_154_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_68_0 dadda_fa_6_68_0/A dadda_fa_6_68_0/B dadda_fa_6_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_69_0/B dadda_fa_7_68_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_71_0 U$$547/Y U$$681/X U$$814/X VGND VGND VPWR VPWR dadda_fa_1_72_6/CIN
+ dadda_fa_1_71_8/A sky130_fd_sc_hd__fa_1
XFILLER_110_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_5_7_1 U$$420/X input234/X VGND VGND VPWR VPWR dadda_fa_6_8_0/B dadda_fa_7_7_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_149_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$360 U$$84/B1 U$$408/A2 U$$634/B1 U$$408/B2 VGND VGND VPWR VPWR U$$361/A sky130_fd_sc_hd__a22o_1
XU$$371 U$$371/A U$$383/B VGND VGND VPWR VPWR U$$371/X sky130_fd_sc_hd__xor2_1
X_629_ _634_/CLK _629_/D VGND VGND VPWR VPWR _629_/Q sky130_fd_sc_hd__dfxtp_4
XU$$382 U$$517/B1 U$$384/A2 U$$382/B1 U$$384/B2 VGND VGND VPWR VPWR U$$383/A sky130_fd_sc_hd__a22o_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$393 U$$393/A U$$393/B VGND VGND VPWR VPWR U$$393/X sky130_fd_sc_hd__xor2_1
XFILLER_199_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_93_1 U$$3252/X U$$3385/X U$$3518/X VGND VGND VPWR VPWR dadda_fa_3_94_0/CIN
+ dadda_fa_3_93_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_195_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_70_0 dadda_fa_5_70_0/A dadda_fa_5_70_0/B dadda_fa_5_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_71_0/A dadda_fa_6_70_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_86_0 U$$3770/X U$$3903/X U$$4036/X VGND VGND VPWR VPWR dadda_fa_3_87_0/B
+ dadda_fa_3_86_2/B sky130_fd_sc_hd__fa_1
Xrepeater1260 U$$4502/A1 VGND VGND VPWR VPWR U$$940/A1 sky130_fd_sc_hd__buf_6
Xrepeater1271 _606_/Q VGND VGND VPWR VPWR U$$3404/A1 sky130_fd_sc_hd__buf_4
Xrepeater1282 U$$3124/B1 VGND VGND VPWR VPWR U$$384/B1 sky130_fd_sc_hd__buf_8
XFILLER_113_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1293 _603_/Q VGND VGND VPWR VPWR U$$2848/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_141_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_49_7 U$$2898/X U$$3031/X VGND VGND VPWR VPWR dadda_fa_2_50_3/A dadda_fa_3_49_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_86_115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_62_7 dadda_fa_1_62_7/A dadda_fa_1_62_7/B dadda_fa_1_62_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_2/CIN dadda_fa_2_62_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_55_6 U$$3176/X U$$3309/X U$$3442/X VGND VGND VPWR VPWR dadda_fa_2_56_2/B
+ dadda_fa_2_55_5/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_48_5 U$$2098/X U$$2231/X U$$2364/X VGND VGND VPWR VPWR dadda_fa_2_49_2/CIN
+ dadda_fa_2_48_5/B sky130_fd_sc_hd__fa_1
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_7_0 dadda_fa_7_7_0/A dadda_fa_7_7_0/B dadda_fa_7_7_0/CIN VGND VGND VPWR
+ VPWR _432_/D _303_/D sky130_fd_sc_hd__fa_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_85_0 dadda_fa_7_85_0/A dadda_fa_7_85_0/B dadda_fa_7_85_0/CIN VGND VGND
+ VPWR VPWR _510_/D _381_/D sky130_fd_sc_hd__fa_1
XFILLER_12_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4108 U$$4108/A U$$4109/A VGND VGND VPWR VPWR U$$4108/X sky130_fd_sc_hd__xor2_1
XU$$4119 U$$4119/A U$$4141/B VGND VGND VPWR VPWR U$$4119/X sky130_fd_sc_hd__xor2_1
XFILLER_150_1242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3407 U$$3407/A U$$3407/B VGND VGND VPWR VPWR U$$3407/X sky130_fd_sc_hd__xor2_1
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3418 U$$3418/A1 U$$3418/A2 U$$4105/A1 U$$3418/B2 VGND VGND VPWR VPWR U$$3419/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_100_0 dadda_fa_6_100_0/A dadda_fa_6_100_0/B dadda_fa_6_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_101_0/B dadda_fa_7_100_0/CIN sky130_fd_sc_hd__fa_1
XU$$3429 U$$3427/Y _666_/Q U$$3425/A U$$3428/X U$$3425/Y VGND VGND VPWR VPWR U$$3429/X
+ sky130_fd_sc_hd__a32o_4
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2706 U$$2706/A U$$2706/B VGND VGND VPWR VPWR U$$2706/X sky130_fd_sc_hd__xor2_1
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2717 U$$2717/A1 U$$2733/A2 U$$3404/A1 U$$2733/B2 VGND VGND VPWR VPWR U$$2718/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2728 U$$2728/A U$$2730/B VGND VGND VPWR VPWR U$$2728/X sky130_fd_sc_hd__xor2_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2739 U$$2739/A VGND VGND VPWR VPWR U$$2739/Y sky130_fd_sc_hd__inv_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ _542_/CLK _414_/D VGND VGND VPWR VPWR _414_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ _476_/CLK _345_/D VGND VGND VPWR VPWR _345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1098 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_498 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_276_ _521_/CLK _276_/D VGND VGND VPWR VPWR _276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_65_5 dadda_fa_2_65_5/A dadda_fa_2_65_5/B dadda_fa_2_65_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_2/A dadda_fa_4_65_0/A sky130_fd_sc_hd__fa_1
XFILLER_151_1039 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater905 U$$4382/B VGND VGND VPWR VPWR U$$4384/A sky130_fd_sc_hd__buf_4
Xrepeater916 U$$4247/A VGND VGND VPWR VPWR U$$4246/A sky130_fd_sc_hd__buf_6
XFILLER_84_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater927 U$$4070/B VGND VGND VPWR VPWR U$$4058/B sky130_fd_sc_hd__buf_6
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater938 _673_/Q VGND VGND VPWR VPWR U$$3943/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_58_4 dadda_fa_2_58_4/A dadda_fa_2_58_4/B dadda_fa_2_58_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/CIN dadda_fa_3_58_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater949 U$$3675/B VGND VGND VPWR VPWR U$$3609/B sky130_fd_sc_hd__buf_6
XU$$3930 _595_/Q U$$3840/X _596_/Q U$$3841/X VGND VGND VPWR VPWR U$$3931/A sky130_fd_sc_hd__a22o_1
XFILLER_25_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3941 U$$3941/A U$$3943/B VGND VGND VPWR VPWR U$$3941/X sky130_fd_sc_hd__xor2_1
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3952 U$$4087/B1 U$$3968/A2 U$$3952/B1 U$$3968/B2 VGND VGND VPWR VPWR U$$3953/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3963 U$$3963/A U$$3965/B VGND VGND VPWR VPWR U$$3963/X sky130_fd_sc_hd__xor2_1
XU$$3974 _674_/Q VGND VGND VPWR VPWR U$$3976/B sky130_fd_sc_hd__inv_1
XU$$3985 U$$4396/A1 U$$4005/A2 U$$4259/B1 U$$4005/B2 VGND VGND VPWR VPWR U$$3986/A
+ sky130_fd_sc_hd__a22o_1
XU$$3996 U$$3996/A U$$4096/B VGND VGND VPWR VPWR U$$3996/X sky130_fd_sc_hd__xor2_1
XFILLER_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_398 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$190 U$$190/A U$$190/B VGND VGND VPWR VPWR U$$190/X sky130_fd_sc_hd__xor2_1
XFILLER_127_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$819_1844 VGND VGND VPWR VPWR U$$819_1844/HI U$$819/B1 sky130_fd_sc_hd__conb_1
XFILLER_119_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_952 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput265 _275_/Q VGND VGND VPWR VPWR o[107] sky130_fd_sc_hd__buf_2
XFILLER_114_551 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput276 _285_/Q VGND VGND VPWR VPWR o[117] sky130_fd_sc_hd__buf_2
XFILLER_47_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1090 U$$1636/B VGND VGND VPWR VPWR U$$1588/B sky130_fd_sc_hd__buf_8
Xoutput287 _295_/Q VGND VGND VPWR VPWR o[127] sky130_fd_sc_hd__buf_2
Xoutput298 _189_/Q VGND VGND VPWR VPWR o[21] sky130_fd_sc_hd__buf_2
XFILLER_141_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_60_4 U$$3585/X U$$3718/X U$$3851/X VGND VGND VPWR VPWR dadda_fa_2_61_1/CIN
+ dadda_fa_2_60_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_53_3 U$$1576/X U$$1709/X U$$1842/X VGND VGND VPWR VPWR dadda_fa_2_54_1/B
+ dadda_fa_2_53_4/B sky130_fd_sc_hd__fa_1
XFILLER_67_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_30_2 dadda_fa_4_30_2/A dadda_fa_4_30_2/B dadda_fa_4_30_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/CIN dadda_fa_5_30_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_46_2 U$$897/X U$$1030/X U$$1163/X VGND VGND VPWR VPWR dadda_fa_2_47_2/B
+ dadda_fa_2_46_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_43_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_23_1 dadda_fa_4_23_1/A dadda_fa_4_23_1/B dadda_fa_4_23_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/B dadda_fa_5_23_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_39_1 U$$484/X U$$617/X U$$750/X VGND VGND VPWR VPWR dadda_fa_2_40_4/B
+ dadda_fa_2_39_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_71_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_16_0 U$$704/X U$$837/X U$$970/X VGND VGND VPWR VPWR dadda_fa_5_17_0/A
+ dadda_fa_5_16_1/A sky130_fd_sc_hd__fa_1
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_582 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_68_3 dadda_fa_3_68_3/A dadda_fa_3_68_3/B dadda_fa_3_68_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_1/B dadda_fa_4_68_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_61_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3204 U$$3204/A U$$3286/B VGND VGND VPWR VPWR U$$3204/X sky130_fd_sc_hd__xor2_1
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3215 U$$3352/A1 U$$3215/A2 U$$3217/A1 U$$3215/B2 VGND VGND VPWR VPWR U$$3216/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3226 U$$3226/A U$$3256/B VGND VGND VPWR VPWR U$$3226/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_85_clk _628_/CLK VGND VGND VPWR VPWR _627_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$19 _443_/Q _315_/Q VGND VGND VPWR VPWR final_adder.U$$147/B1 final_adder.U$$641/A
+ sky130_fd_sc_hd__ha_2
XU$$3237 U$$3374/A1 U$$3285/A2 U$$4472/A1 U$$3285/B2 VGND VGND VPWR VPWR U$$3238/A
+ sky130_fd_sc_hd__a22o_1
XU$$2503 U$$2503/A U$$2551/B VGND VGND VPWR VPWR U$$2503/X sky130_fd_sc_hd__xor2_1
XU$$3248 U$$3248/A U$$3256/B VGND VGND VPWR VPWR U$$3248/X sky130_fd_sc_hd__xor2_1
XU$$3259 _602_/Q U$$3263/A2 _603_/Q U$$3263/B2 VGND VGND VPWR VPWR U$$3260/A sky130_fd_sc_hd__a22o_1
XFILLER_46_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2514 U$$2786/B1 U$$2516/A2 U$$3475/A1 U$$2516/B2 VGND VGND VPWR VPWR U$$2515/A
+ sky130_fd_sc_hd__a22o_1
XU$$2525 U$$2525/A U$$2531/B VGND VGND VPWR VPWR U$$2525/X sky130_fd_sc_hd__xor2_1
XU$$2536 U$$3769/A1 U$$2470/X U$$3769/B1 U$$2471/X VGND VGND VPWR VPWR U$$2537/A sky130_fd_sc_hd__a22o_1
XFILLER_74_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1802 U$$1802/A U$$1852/B VGND VGND VPWR VPWR U$$1802/X sky130_fd_sc_hd__xor2_1
XU$$2547 U$$2547/A U$$2551/B VGND VGND VPWR VPWR U$$2547/X sky130_fd_sc_hd__xor2_1
XFILLER_62_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1813 U$$715/B1 U$$1855/A2 U$$582/A1 U$$1855/B2 VGND VGND VPWR VPWR U$$1814/A sky130_fd_sc_hd__a22o_1
XU$$2558 U$$3789/B1 U$$2588/A2 U$$916/A1 U$$2588/B2 VGND VGND VPWR VPWR U$$2559/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1824 U$$1824/A U$$1874/B VGND VGND VPWR VPWR U$$1824/X sky130_fd_sc_hd__xor2_1
XU$$2569 U$$2569/A U$$2583/B VGND VGND VPWR VPWR U$$2569/X sky130_fd_sc_hd__xor2_1
XU$$1835 U$$3342/A1 U$$1843/A2 U$$467/A1 U$$1843/B2 VGND VGND VPWR VPWR U$$1836/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1846 U$$1846/A U$$1917/A VGND VGND VPWR VPWR U$$1846/X sky130_fd_sc_hd__xor2_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1857 U$$624/A1 U$$1785/X U$$624/B1 U$$1786/X VGND VGND VPWR VPWR U$$1858/A sky130_fd_sc_hd__a22o_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1868 U$$1868/A U$$1870/B VGND VGND VPWR VPWR U$$1868/X sky130_fd_sc_hd__xor2_1
XFILLER_15_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1879 U$$3112/A1 U$$1907/A2 U$$922/A1 U$$1907/B2 VGND VGND VPWR VPWR U$$1880/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_328_ _478_/CLK _328_/D VGND VGND VPWR VPWR _328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_259_ _379_/CLK _259_/D VGND VGND VPWR VPWR _259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_70_3 dadda_fa_2_70_3/A dadda_fa_2_70_3/B dadda_fa_2_70_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/B dadda_fa_3_70_3/B sky130_fd_sc_hd__fa_1
Xdadda_fa_2_63_2 dadda_fa_2_63_2/A dadda_fa_2_63_2/B dadda_fa_2_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/A dadda_fa_3_63_3/A sky130_fd_sc_hd__fa_1
XFILLER_69_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater702 U$$3978/X VGND VGND VPWR VPWR U$$4071/B2 sky130_fd_sc_hd__buf_6
Xrepeater713 U$$3795/B2 VGND VGND VPWR VPWR U$$3785/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$509 final_adder.U$$636/A final_adder.U$$636/B final_adder.U$$509/B1
+ VGND VGND VPWR VPWR final_adder.U$$637/B sky130_fd_sc_hd__a21o_1
XFILLER_96_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater724 U$$3567/X VGND VGND VPWR VPWR U$$3664/B2 sky130_fd_sc_hd__buf_4
XFILLER_84_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_40_1 dadda_fa_5_40_1/A dadda_fa_5_40_1/B dadda_fa_5_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_41_0/B dadda_fa_7_40_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_56_1 dadda_fa_2_56_1/A dadda_fa_2_56_1/B dadda_fa_2_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_0/CIN dadda_fa_3_56_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater735 U$$3293/X VGND VGND VPWR VPWR U$$3418/B2 sky130_fd_sc_hd__buf_6
Xrepeater746 U$$3283/B2 VGND VGND VPWR VPWR U$$3285/B2 sky130_fd_sc_hd__buf_6
XFILLER_38_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater757 U$$3148/B2 VGND VGND VPWR VPWR U$$3144/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_33_0 dadda_fa_5_33_0/A dadda_fa_5_33_0/B dadda_fa_5_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_34_0/A dadda_fa_6_33_0/CIN sky130_fd_sc_hd__fa_2
XU$$4450 U$$4450/A1 U$$4388/X U$$4450/B1 U$$4454/B2 VGND VGND VPWR VPWR U$$4451/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater768 U$$334/B2 VGND VGND VPWR VPWR U$$308/B2 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_76_clk _628_/CLK VGND VGND VPWR VPWR _679_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$4461 U$$4461/A U$$4461/B VGND VGND VPWR VPWR U$$4461/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_49_0 U$$3164/X U$$3297/X input200/X VGND VGND VPWR VPWR dadda_fa_3_50_0/B
+ dadda_fa_3_49_2/B sky130_fd_sc_hd__fa_1
Xrepeater779 U$$2745/X VGND VGND VPWR VPWR U$$2832/B2 sky130_fd_sc_hd__buf_6
XFILLER_49_192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4472 U$$4472/A1 U$$4388/X U$$4472/B1 U$$4480/B2 VGND VGND VPWR VPWR U$$4473/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4483 U$$4483/A U$$4483/B VGND VGND VPWR VPWR U$$4483/X sky130_fd_sc_hd__xor2_1
XU$$4494 U$$932/A1 U$$4388/X U$$4494/B1 U$$4496/B2 VGND VGND VPWR VPWR U$$4495/A sky130_fd_sc_hd__a22o_1
XU$$3760 U$$3760/A U$$3760/B VGND VGND VPWR VPWR U$$3760/X sky130_fd_sc_hd__xor2_1
XU$$3771 U$$4045/A1 U$$3823/A2 U$$3771/B1 U$$3823/B2 VGND VGND VPWR VPWR U$$3772/A
+ sky130_fd_sc_hd__a22o_1
XU$$3782 U$$3782/A U$$3800/B VGND VGND VPWR VPWR U$$3782/X sky130_fd_sc_hd__xor2_1
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3793 _595_/Q U$$3795/A2 _596_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3794/A sky130_fd_sc_hd__a22o_1
XFILLER_197_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_78_2 dadda_fa_4_78_2/A dadda_fa_4_78_2/B dadda_fa_4_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/CIN dadda_fa_5_78_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_48_0 dadda_fa_7_48_0/A dadda_fa_7_48_0/B dadda_fa_7_48_0/CIN VGND VGND
+ VPWR VPWR _473_/D _344_/D sky130_fd_sc_hd__fa_2
XFILLER_48_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_51_0 U$$109/X U$$242/X U$$375/X VGND VGND VPWR VPWR dadda_fa_2_52_0/B
+ dadda_fa_2_51_3/B sky130_fd_sc_hd__fa_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_clk _369_/CLK VGND VGND VPWR VPWR _558_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$904 U$$80/B1 U$$906/A2 U$$906/A1 U$$906/B2 VGND VGND VPWR VPWR U$$905/A sky130_fd_sc_hd__a22o_1
XFILLER_28_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$915 U$$915/A U$$958/A VGND VGND VPWR VPWR U$$915/X sky130_fd_sc_hd__xor2_1
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$926 U$$926/A1 U$$928/A2 U$$928/A1 U$$928/B2 VGND VGND VPWR VPWR U$$927/A sky130_fd_sc_hd__a22o_1
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$937 U$$937/A _629_/Q VGND VGND VPWR VPWR U$$937/X sky130_fd_sc_hd__xor2_1
XU$$948 U$$948/A1 U$$948/A2 U$$948/B1 U$$948/B2 VGND VGND VPWR VPWR U$$949/A sky130_fd_sc_hd__a22o_1
XFILLER_28_387 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$959 _629_/Q VGND VGND VPWR VPWR U$$959/Y sky130_fd_sc_hd__inv_1
XU$$1109 U$$1109/A U$$1151/B VGND VGND VPWR VPWR U$$1109/X sky130_fd_sc_hd__xor2_1
XFILLER_203_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1076 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_80_2 dadda_fa_3_80_2/A dadda_fa_3_80_2/B dadda_fa_3_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_1/A dadda_fa_4_80_2/B sky130_fd_sc_hd__fa_1
XFILLER_30_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_73_1 dadda_fa_3_73_1/A dadda_fa_3_73_1/B dadda_fa_3_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_0/CIN dadda_fa_4_73_2/A sky130_fd_sc_hd__fa_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_50_0 dadda_fa_6_50_0/A dadda_fa_6_50_0/B dadda_fa_6_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_51_0/B dadda_fa_7_50_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_66_0 dadda_fa_3_66_0/A dadda_fa_3_66_0/B dadda_fa_3_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_0/B dadda_fa_4_66_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3001 U$$3412/A1 U$$3005/A2 U$$3412/B1 U$$3005/B2 VGND VGND VPWR VPWR U$$3002/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3012 U$$3012/A _659_/Q VGND VGND VPWR VPWR U$$3012/X sky130_fd_sc_hd__xor2_1
XU$$3023 U$$3023/A U$$3065/B VGND VGND VPWR VPWR U$$3023/X sky130_fd_sc_hd__xor2_1
XU$$3034 U$$3445/A1 U$$3046/A2 U$$3310/A1 U$$3046/B2 VGND VGND VPWR VPWR U$$3035/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3045 U$$3045/A U$$3083/B VGND VGND VPWR VPWR U$$3045/X sky130_fd_sc_hd__xor2_1
XFILLER_75_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2300 U$$2983/B1 U$$2302/A2 U$$2848/B1 U$$2302/B2 VGND VGND VPWR VPWR U$$2301/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3056 U$$3193/A1 U$$3066/A2 U$$3056/B1 U$$3066/B2 VGND VGND VPWR VPWR U$$3057/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2311 U$$2311/A U$$2321/B VGND VGND VPWR VPWR U$$2311/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_102_1 dadda_fa_4_102_1/A dadda_fa_4_102_1/B dadda_fa_4_102_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/B dadda_fa_5_102_1/B sky130_fd_sc_hd__fa_1
XFILLER_207_466 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2322 U$$2459/A1 U$$2326/A2 U$$2459/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2323/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3067 U$$3067/A U$$3107/B VGND VGND VPWR VPWR U$$3067/X sky130_fd_sc_hd__xor2_1
XU$$2333 U$$2331/Y _650_/Q _649_/Q U$$2332/X U$$2329/Y VGND VGND VPWR VPWR U$$2333/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3078 U$$4448/A1 U$$3082/A2 U$$3626/B1 U$$3082/B2 VGND VGND VPWR VPWR U$$3079/A
+ sky130_fd_sc_hd__a22o_1
XU$$3089 U$$3089/A U$$3121/B VGND VGND VPWR VPWR U$$3089/X sky130_fd_sc_hd__xor2_1
XU$$2344 U$$2344/A U$$2366/B VGND VGND VPWR VPWR U$$2344/X sky130_fd_sc_hd__xor2_1
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2355 U$$3451/A1 U$$2395/A2 U$$3453/A1 U$$2395/B2 VGND VGND VPWR VPWR U$$2356/A
+ sky130_fd_sc_hd__a22o_1
XU$$1610 U$$1610/A U$$1636/B VGND VGND VPWR VPWR U$$1610/X sky130_fd_sc_hd__xor2_1
XU$$1621 U$$2991/A1 U$$1627/A2 U$$251/B1 U$$1627/B2 VGND VGND VPWR VPWR U$$1622/A
+ sky130_fd_sc_hd__a22o_1
XU$$2366 U$$2366/A U$$2366/B VGND VGND VPWR VPWR U$$2366/X sky130_fd_sc_hd__xor2_1
XFILLER_62_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1632 U$$1632/A U$$1636/B VGND VGND VPWR VPWR U$$1632/X sky130_fd_sc_hd__xor2_1
XFILLER_62_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2377 U$$4156/B1 U$$2423/A2 U$$3884/B1 U$$2423/B2 VGND VGND VPWR VPWR U$$2378/A
+ sky130_fd_sc_hd__a22o_1
XU$$1643 _639_/Q VGND VGND VPWR VPWR U$$1643/Y sky130_fd_sc_hd__inv_1
XFILLER_62_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2388 U$$2388/A U$$2388/B VGND VGND VPWR VPWR U$$2388/X sky130_fd_sc_hd__xor2_1
XU$$2399 U$$890/B1 U$$2437/A2 U$$757/A1 U$$2437/B2 VGND VGND VPWR VPWR U$$2400/A sky130_fd_sc_hd__a22o_1
XU$$1654 U$$695/A1 U$$1684/A2 U$$2613/B1 U$$1684/B2 VGND VGND VPWR VPWR U$$1655/A
+ sky130_fd_sc_hd__a22o_1
XU$$1665 U$$1665/A U$$1687/B VGND VGND VPWR VPWR U$$1665/X sky130_fd_sc_hd__xor2_1
XU$$1676 U$$715/B1 U$$1718/A2 U$$582/A1 U$$1718/B2 VGND VGND VPWR VPWR U$$1677/A sky130_fd_sc_hd__a22o_1
XFILLER_163_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1687 U$$1687/A U$$1687/B VGND VGND VPWR VPWR U$$1687/X sky130_fd_sc_hd__xor2_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_123_0 dadda_fa_7_123_0/A dadda_fa_7_123_0/B dadda_fa_7_123_0/CIN VGND
+ VGND VPWR VPWR _548_/D _419_/D sky130_fd_sc_hd__fa_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1698 U$$3342/A1 U$$1718/A2 U$$467/A1 U$$1718/B2 VGND VGND VPWR VPWR U$$1699/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_88_1 dadda_fa_5_88_1/A dadda_fa_5_88_1/B dadda_fa_5_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_89_0/B dadda_fa_7_88_0/A sky130_fd_sc_hd__fa_1
XFILLER_116_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$306 final_adder.U$$306/A final_adder.U$$306/B VGND VGND VPWR VPWR
+ final_adder.U$$344/A sky130_fd_sc_hd__and2_1
XFILLER_131_1218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater510 U$$3018/X VGND VGND VPWR VPWR U$$3148/A2 sky130_fd_sc_hd__buf_4
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$317 final_adder.U$$316/A final_adder.U$$249/X final_adder.U$$251/X
+ VGND VGND VPWR VPWR final_adder.U$$317/X sky130_fd_sc_hd__a21o_1
Xrepeater521 U$$398/A2 VGND VGND VPWR VPWR U$$334/A2 sky130_fd_sc_hd__buf_6
XFILLER_69_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$328 final_adder.U$$328/A final_adder.U$$328/B VGND VGND VPWR VPWR
+ final_adder.U$$356/B sky130_fd_sc_hd__and2_1
Xrepeater532 U$$2866/A2 VGND VGND VPWR VPWR U$$2856/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$339 final_adder.U$$338/A final_adder.U$$293/X final_adder.U$$295/X
+ VGND VGND VPWR VPWR final_adder.U$$339/X sky130_fd_sc_hd__a21o_1
Xrepeater543 U$$2566/A2 VGND VGND VPWR VPWR U$$2550/A2 sky130_fd_sc_hd__buf_4
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_49_clk _369_/CLK VGND VGND VPWR VPWR _519_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater554 U$$2437/A2 VGND VGND VPWR VPWR U$$2395/A2 sky130_fd_sc_hd__buf_4
XFILLER_211_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater565 U$$2318/A2 VGND VGND VPWR VPWR U$$2326/A2 sky130_fd_sc_hd__buf_4
XFILLER_38_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater576 U$$1982/A2 VGND VGND VPWR VPWR U$$1976/A2 sky130_fd_sc_hd__buf_4
Xrepeater587 U$$1915/A2 VGND VGND VPWR VPWR U$$1897/A2 sky130_fd_sc_hd__buf_6
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4280 U$$4280/A U$$4322/B VGND VGND VPWR VPWR U$$4280/X sky130_fd_sc_hd__xor2_1
Xrepeater598 U$$1648/X VGND VGND VPWR VPWR U$$1778/A2 sky130_fd_sc_hd__buf_6
XFILLER_38_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_482 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4291 U$$4291/A1 U$$4311/A2 U$$4293/A1 U$$4311/B2 VGND VGND VPWR VPWR U$$4292/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3590 U$$4136/B1 U$$3636/A2 U$$4003/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3591/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_833 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_90_1 dadda_fa_4_90_1/A dadda_fa_4_90_1/B dadda_fa_4_90_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/B dadda_fa_5_90_1/B sky130_fd_sc_hd__fa_1
XFILLER_107_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_83_0 dadda_fa_4_83_0/A dadda_fa_4_83_0/B dadda_fa_4_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/A dadda_fa_5_83_1/A sky130_fd_sc_hd__fa_1
XFILLER_162_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_104_3 dadda_fa_3_104_3/A dadda_fa_3_104_3/B dadda_fa_3_104_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_105_1/B dadda_fa_4_104_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$701 U$$838/A1 U$$725/A2 U$$840/A1 U$$725/B2 VGND VGND VPWR VPWR U$$702/A sky130_fd_sc_hd__a22o_1
XFILLER_57_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_662_ _662_/CLK _662_/D VGND VGND VPWR VPWR _662_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$712 U$$712/A U$$766/B VGND VGND VPWR VPWR U$$712/X sky130_fd_sc_hd__xor2_1
XU$$723 U$$38/A1 U$$725/A2 U$$40/A1 U$$725/B2 VGND VGND VPWR VPWR U$$724/A sky130_fd_sc_hd__a22o_1
XFILLER_57_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$734 U$$734/A U$$760/B VGND VGND VPWR VPWR U$$734/X sky130_fd_sc_hd__xor2_1
XU$$745 U$$745/A1 U$$747/A2 U$$882/B1 U$$747/B2 VGND VGND VPWR VPWR U$$746/A sky130_fd_sc_hd__a22o_1
XFILLER_112_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_593_ _596_/CLK _593_/D VGND VGND VPWR VPWR _593_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$756 U$$756/A U$$796/B VGND VGND VPWR VPWR U$$756/X sky130_fd_sc_hd__xor2_1
XFILLER_45_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$767 U$$82/A1 U$$783/A2 U$$84/A1 U$$783/B2 VGND VGND VPWR VPWR U$$768/A sky130_fd_sc_hd__a22o_1
XU$$778 U$$778/A U$$816/B VGND VGND VPWR VPWR U$$778/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$789 U$$924/B1 U$$809/A2 U$$791/A1 U$$809/B2 VGND VGND VPWR VPWR U$$790/A sky130_fd_sc_hd__a22o_1
XFILLER_189_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_98_0 dadda_fa_6_98_0/A dadda_fa_6_98_0/B dadda_fa_6_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_99_0/B dadda_fa_7_98_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_145_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1601 U$$3046/B1 VGND VGND VPWR VPWR U$$4418/A1 sky130_fd_sc_hd__buf_6
XFILLER_144_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_6 _456_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1612 U$$4140/A1 VGND VGND VPWR VPWR U$$715/A1 sky130_fd_sc_hd__buf_6
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1623 U$$3453/A1 VGND VGND VPWR VPWR U$$987/A1 sky130_fd_sc_hd__buf_6
Xrepeater1634 U$$4273/A1 VGND VGND VPWR VPWR U$$3312/B1 sky130_fd_sc_hd__buf_8
Xrepeater1645 _560_/Q VGND VGND VPWR VPWR U$$3447/B1 sky130_fd_sc_hd__buf_8
XFILLER_152_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1656 U$$3717/B1 VGND VGND VPWR VPWR U$$429/B1 sky130_fd_sc_hd__buf_4
Xrepeater1667 U$$2893/B1 VGND VGND VPWR VPWR U$$2895/A1 sky130_fd_sc_hd__buf_6
XFILLER_193_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1678 _556_/Q VGND VGND VPWR VPWR U$$3713/B1 sky130_fd_sc_hd__buf_8
Xrepeater1689 U$$3024/B1 VGND VGND VPWR VPWR U$$971/A1 sky130_fd_sc_hd__buf_4
XFILLER_113_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1040 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_40_4 dadda_fa_2_40_4/A dadda_fa_2_40_4/B dadda_fa_2_40_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_41_1/CIN dadda_fa_3_40_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4463_1810 VGND VGND VPWR VPWR U$$4463_1810/HI U$$4463/B sky130_fd_sc_hd__conb_1
Xdadda_fa_2_33_3 U$$1270/X U$$1403/X U$$1536/X VGND VGND VPWR VPWR dadda_fa_3_34_1/B
+ dadda_fa_3_33_3/B sky130_fd_sc_hd__fa_1
XFILLER_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2130 U$$2130/A U$$2130/B VGND VGND VPWR VPWR U$$2130/X sky130_fd_sc_hd__xor2_1
XFILLER_63_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2141 U$$3783/B1 U$$2169/A2 U$$2963/B1 U$$2169/B2 VGND VGND VPWR VPWR U$$2142/A
+ sky130_fd_sc_hd__a22o_1
XU$$2152 U$$2152/A U$$2191/A VGND VGND VPWR VPWR U$$2152/X sky130_fd_sc_hd__xor2_1
XU$$2163 U$$2983/B1 U$$2189/A2 U$$2848/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2164/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2174 U$$2174/A U$$2174/B VGND VGND VPWR VPWR U$$2174/X sky130_fd_sc_hd__xor2_1
XU$$1440 U$$344/A1 U$$1442/A2 U$$3221/B1 U$$1442/B2 VGND VGND VPWR VPWR U$$1441/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2185 U$$952/A1 U$$2185/A2 U$$2459/B1 U$$2185/B2 VGND VGND VPWR VPWR U$$2186/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1451 U$$1451/A U$$1479/B VGND VGND VPWR VPWR U$$1451/X sky130_fd_sc_hd__xor2_1
XU$$2196 U$$2194/Y _648_/Q _647_/Q U$$2195/X U$$2192/Y VGND VGND VPWR VPWR U$$2196/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_204_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1462 U$$92/A1 U$$1474/A2 U$$94/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1463/A sky130_fd_sc_hd__a22o_1
XU$$1473 U$$1473/A U$$1475/B VGND VGND VPWR VPWR U$$1473/X sky130_fd_sc_hd__xor2_1
XFILLER_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1484 U$$251/A1 U$$1486/A2 U$$251/B1 U$$1486/B2 VGND VGND VPWR VPWR U$$1485/A sky130_fd_sc_hd__a22o_1
XU$$1495 U$$1495/A U$$1501/B VGND VGND VPWR VPWR U$$1495/X sky130_fd_sc_hd__xor2_1
XFILLER_187_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_78_5 U$$3222/X U$$3355/X U$$3488/X VGND VGND VPWR VPWR dadda_fa_2_79_2/A
+ dadda_fa_2_78_5/A sky130_fd_sc_hd__fa_1
XFILLER_170_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$103 _527_/Q _399_/Q VGND VGND VPWR VPWR final_adder.U$$231/B1 final_adder.U$$725/A
+ sky130_fd_sc_hd__ha_1
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$114 _538_/Q _410_/Q VGND VGND VPWR VPWR final_adder.U$$609/B1 final_adder.U$$736/A
+ sky130_fd_sc_hd__ha_2
XFILLER_44_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$125 _549_/Q _421_/Q VGND VGND VPWR VPWR final_adder.U$$253/B1 final_adder.U$$747/A
+ sky130_fd_sc_hd__ha_2
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$136 final_adder.U$$9/SUM final_adder.U$$8/SUM VGND VGND VPWR VPWR
+ final_adder.U$$260/B sky130_fd_sc_hd__and2_1
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$147 final_adder.U$$641/A final_adder.U$$513/B1 final_adder.U$$147/B1
+ VGND VGND VPWR VPWR final_adder.U$$147/X sky130_fd_sc_hd__a21o_1
XFILLER_79_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$158 final_adder.U$$653/A final_adder.U$$652/A VGND VGND VPWR VPWR
+ final_adder.U$$270/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$169 final_adder.U$$663/A final_adder.U$$535/B1 final_adder.U$$169/B1
+ VGND VGND VPWR VPWR final_adder.U$$169/X sky130_fd_sc_hd__a21o_1
XFILLER_39_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater395 U$$896/A2 VGND VGND VPWR VPWR U$$878/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_282 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_579 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_76 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_102_0 U$$4068/X U$$4201/X U$$4334/X VGND VGND VPWR VPWR dadda_fa_4_103_0/B
+ dadda_fa_4_102_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_891 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput110 b[50] VGND VGND VPWR VPWR _602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput121 b[60] VGND VGND VPWR VPWR _612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput132 c[102] VGND VGND VPWR VPWR input132/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_50_3 dadda_fa_3_50_3/A dadda_fa_3_50_3/B dadda_fa_3_50_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_1/B dadda_fa_4_50_2/CIN sky130_fd_sc_hd__fa_1
Xinput143 c[112] VGND VGND VPWR VPWR input143/X sky130_fd_sc_hd__clkbuf_1
XTAP_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_66_3 U$$1336/X U$$1469/X U$$1602/X VGND VGND VPWR VPWR dadda_fa_1_67_6/B
+ dadda_fa_1_66_8/B sky130_fd_sc_hd__fa_1
Xinput154 c[122] VGND VGND VPWR VPWR input154/X sky130_fd_sc_hd__clkbuf_1
XTAP_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput165 c[17] VGND VGND VPWR VPWR input165/X sky130_fd_sc_hd__clkbuf_1
XTAP_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput176 c[27] VGND VGND VPWR VPWR input176/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_3_43_2 dadda_fa_3_43_2/A dadda_fa_3_43_2/B dadda_fa_3_43_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_1/A dadda_fa_4_43_2/B sky130_fd_sc_hd__fa_1
XTAP_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput187 c[37] VGND VGND VPWR VPWR input187/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput198 c[47] VGND VGND VPWR VPWR input198/X sky130_fd_sc_hd__buf_2
XFILLER_64_728 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_59_2 U$$923/X U$$1056/X U$$1189/X VGND VGND VPWR VPWR dadda_fa_1_60_7/A
+ dadda_fa_1_59_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$670 final_adder.U$$670/A final_adder.U$$670/B VGND VGND VPWR VPWR
+ _216_/D sky130_fd_sc_hd__xor2_1
XTAP_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$681 final_adder.U$$681/A final_adder.U$$681/B VGND VGND VPWR VPWR
+ _227_/D sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_36_1 dadda_fa_3_36_1/A dadda_fa_3_36_1/B dadda_fa_3_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_0/CIN dadda_fa_4_36_2/A sky130_fd_sc_hd__fa_1
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$520 U$$520/A U$$547/A VGND VGND VPWR VPWR U$$520/X sky130_fd_sc_hd__xor2_1
XTAP_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_645_ _648_/CLK _645_/D VGND VGND VPWR VPWR _645_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$531 U$$805/A1 U$$415/X U$$805/B1 U$$416/X VGND VGND VPWR VPWR U$$532/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$692 final_adder.U$$692/A final_adder.U$$692/B VGND VGND VPWR VPWR
+ _238_/D sky130_fd_sc_hd__xor2_4
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$542 U$$542/A U$$547/A VGND VGND VPWR VPWR U$$542/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_13_0 dadda_fa_6_13_0/A dadda_fa_6_13_0/B dadda_fa_6_13_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_14_0/B dadda_fa_7_13_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$553 U$$551/B _623_/Q _624_/Q U$$548/Y VGND VGND VPWR VPWR U$$553/X sky130_fd_sc_hd__a22o_2
XFILLER_72_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$564 U$$838/A1 U$$574/A2 U$$840/A1 U$$574/B2 VGND VGND VPWR VPWR U$$565/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_29_0 U$$1528/X U$$1661/X U$$1794/X VGND VGND VPWR VPWR dadda_fa_4_30_0/B
+ dadda_fa_4_29_1/CIN sky130_fd_sc_hd__fa_1
XU$$575 U$$575/A U$$589/B VGND VGND VPWR VPWR U$$575/X sky130_fd_sc_hd__xor2_1
X_576_ _582_/CLK _576_/D VGND VGND VPWR VPWR _576_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_186_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$586 U$$997/A1 U$$600/A2 U$$999/A1 U$$600/B2 VGND VGND VPWR VPWR U$$587/A sky130_fd_sc_hd__a22o_1
XU$$597 U$$597/A U$$665/B VGND VGND VPWR VPWR U$$597/X sky130_fd_sc_hd__xor2_1
XFILLER_72_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$956_1846 VGND VGND VPWR VPWR U$$956_1846/HI U$$956/B1 sky130_fd_sc_hd__conb_1
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4493_1825 VGND VGND VPWR VPWR U$$4493_1825/HI U$$4493/B sky130_fd_sc_hd__conb_1
Xdadda_fa_2_95_5 input251/X dadda_fa_2_95_5/B dadda_fa_2_95_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_96_2/A dadda_fa_4_95_0/A sky130_fd_sc_hd__fa_1
XFILLER_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1420 U$$900/A1 VGND VGND VPWR VPWR U$$761/B1 sky130_fd_sc_hd__buf_6
Xrepeater1431 U$$3638/A1 VGND VGND VPWR VPWR U$$624/A1 sky130_fd_sc_hd__buf_4
Xrepeater1442 _585_/Q VGND VGND VPWR VPWR U$$4456/B1 sky130_fd_sc_hd__buf_4
Xrepeater1453 U$$3358/A1 VGND VGND VPWR VPWR U$$3495/A1 sky130_fd_sc_hd__buf_6
XFILLER_114_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1464 _582_/Q VGND VGND VPWR VPWR U$$4450/B1 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_2_88_4 dadda_fa_2_88_4/A dadda_fa_2_88_4/B dadda_fa_2_88_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_1/CIN dadda_fa_3_88_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1475 _580_/Q VGND VGND VPWR VPWR U$$3352/A1 sky130_fd_sc_hd__buf_6
Xrepeater1486 U$$3896/B1 VGND VGND VPWR VPWR U$$334/B1 sky130_fd_sc_hd__buf_6
XFILLER_207_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1497 U$$4444/A1 VGND VGND VPWR VPWR U$$4031/B1 sky130_fd_sc_hd__buf_6
XFILLER_114_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_25_1 U$$456/X U$$589/X VGND VGND VPWR VPWR dadda_fa_3_26_3/A dadda_fa_4_25_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_67_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_31_0 U$$69/X U$$202/X U$$335/X VGND VGND VPWR VPWR dadda_fa_3_32_0/CIN
+ dadda_fa_3_31_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1270 U$$1270/A U$$1280/B VGND VGND VPWR VPWR U$$1270/X sky130_fd_sc_hd__xor2_1
XFILLER_149_811 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1281 U$$4158/A1 U$$1295/A2 U$$50/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1282/A sky130_fd_sc_hd__a22o_1
XFILLER_195_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1292 U$$1292/A U$$1292/B VGND VGND VPWR VPWR U$$1292/X sky130_fd_sc_hd__xor2_1
XFILLER_148_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_118_0 dadda_fa_5_118_0/A dadda_fa_5_118_0/B dadda_fa_5_118_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_119_0/A dadda_fa_6_118_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_699 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_3 U$$2567/X U$$2700/X U$$2833/X VGND VGND VPWR VPWR dadda_fa_2_84_2/CIN
+ dadda_fa_2_83_5/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_60_2 dadda_fa_4_60_2/A dadda_fa_4_60_2/B dadda_fa_4_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/CIN dadda_fa_5_60_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_76_2 U$$2287/X U$$2420/X U$$2553/X VGND VGND VPWR VPWR dadda_fa_2_77_1/A
+ dadda_fa_2_76_4/A sky130_fd_sc_hd__fa_1
XFILLER_77_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_53_1 dadda_fa_4_53_1/A dadda_fa_4_53_1/B dadda_fa_4_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/B dadda_fa_5_53_1/B sky130_fd_sc_hd__fa_1
XFILLER_58_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_69_1 U$$2805/X U$$2938/X U$$3071/X VGND VGND VPWR VPWR dadda_fa_2_70_0/CIN
+ dadda_fa_2_69_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_30_0 dadda_fa_7_30_0/A dadda_fa_7_30_0/B dadda_fa_7_30_0/CIN VGND VGND
+ VPWR VPWR _455_/D _326_/D sky130_fd_sc_hd__fa_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_46_0 dadda_fa_4_46_0/A dadda_fa_4_46_0/B dadda_fa_4_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/A dadda_fa_5_46_1/A sky130_fd_sc_hd__fa_1
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _190_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_430_ _431_/CLK _430_/D VGND VGND VPWR VPWR _430_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_248 _194_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_259 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_580 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_361_ _491_/CLK _361_/D VGND VGND VPWR VPWR _361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_292_ _615_/CLK _292_/D VGND VGND VPWR VPWR _292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_98_3 dadda_fa_3_98_3/A dadda_fa_3_98_3/B dadda_fa_3_98_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_1/B dadda_fa_4_98_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_72_3 U$$1747/X U$$1880/X VGND VGND VPWR VPWR dadda_fa_1_73_8/A dadda_fa_2_72_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_71_1 U$$947/X U$$1080/X U$$1213/X VGND VGND VPWR VPWR dadda_fa_1_72_7/A
+ dadda_fa_1_71_8/B sky130_fd_sc_hd__fa_1
XTAP_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_64_0 U$$135/X U$$268/X U$$401/X VGND VGND VPWR VPWR dadda_fa_1_65_5/B
+ dadda_fa_1_64_7/B sky130_fd_sc_hd__fa_1
XTAP_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$350 U$$898/A1 U$$350/A2 U$$900/A1 U$$350/B2 VGND VGND VPWR VPWR U$$351/A sky130_fd_sc_hd__a22o_1
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_628_ _628_/CLK _628_/D VGND VGND VPWR VPWR _628_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$361 U$$361/A U$$410/A VGND VGND VPWR VPWR U$$361/X sky130_fd_sc_hd__xor2_1
XU$$372 U$$781/B1 U$$384/A2 U$$648/A1 U$$384/B2 VGND VGND VPWR VPWR U$$373/A sky130_fd_sc_hd__a22o_1
XU$$383 U$$383/A U$$383/B VGND VGND VPWR VPWR U$$383/X sky130_fd_sc_hd__xor2_1
XU$$394 U$$942/A1 U$$408/A2 U$$942/B1 U$$408/B2 VGND VGND VPWR VPWR U$$395/A sky130_fd_sc_hd__a22o_1
X_559_ _559_/CLK _559_/D VGND VGND VPWR VPWR _559_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_199_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_93_2 U$$3651/X U$$3784/X U$$3917/X VGND VGND VPWR VPWR dadda_fa_3_94_1/A
+ dadda_fa_3_93_3/A sky130_fd_sc_hd__fa_1
Xrepeater1250 U$$4228/B1 VGND VGND VPWR VPWR U$$805/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_70_1 dadda_fa_5_70_1/A dadda_fa_5_70_1/B dadda_fa_5_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_71_0/B dadda_fa_7_70_0/A sky130_fd_sc_hd__fa_1
Xrepeater1261 U$$3132/A1 VGND VGND VPWR VPWR U$$4502/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_86_1 U$$4169/X U$$4302/X U$$4435/X VGND VGND VPWR VPWR dadda_fa_3_87_0/CIN
+ dadda_fa_3_86_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater1272 _606_/Q VGND VGND VPWR VPWR U$$2991/B1 sky130_fd_sc_hd__buf_6
Xrepeater1283 _604_/Q VGND VGND VPWR VPWR U$$3124/B1 sky130_fd_sc_hd__buf_4
Xrepeater1294 U$$4357/A1 VGND VGND VPWR VPWR U$$932/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_63_0 dadda_fa_5_63_0/A dadda_fa_5_63_0/B dadda_fa_5_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_64_0/A dadda_fa_6_63_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_79_0 dadda_fa_2_79_0/A dadda_fa_2_79_0/B dadda_fa_2_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_0/B dadda_fa_3_79_2/B sky130_fd_sc_hd__fa_1
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_8 dadda_fa_1_62_8/A dadda_fa_1_62_8/B dadda_fa_1_62_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_3/A dadda_fa_3_62_0/A sky130_fd_sc_hd__fa_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_812 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_55_7 U$$3575/X U$$3708/X input207/X VGND VGND VPWR VPWR dadda_fa_2_56_2/CIN
+ dadda_fa_2_55_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_48_6 U$$2497/X U$$2630/X U$$2763/X VGND VGND VPWR VPWR dadda_fa_2_49_3/A
+ dadda_fa_2_48_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_167_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_56 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_78_0 dadda_fa_7_78_0/A dadda_fa_7_78_0/B dadda_fa_7_78_0/CIN VGND VGND
+ VPWR VPWR _503_/D _374_/D sky130_fd_sc_hd__fa_1
XFILLER_191_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_81_0 U$$1232/Y U$$1366/X U$$1499/X VGND VGND VPWR VPWR dadda_fa_2_82_1/A
+ dadda_fa_2_81_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_144_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_606 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4109 U$$4109/A VGND VGND VPWR VPWR U$$4109/Y sky130_fd_sc_hd__inv_1
XFILLER_63_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3408 U$$4504/A1 U$$3408/A2 U$$4506/A1 U$$3408/B2 VGND VGND VPWR VPWR U$$3409/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3419 U$$3419/A U$$3424/A VGND VGND VPWR VPWR U$$3419/X sky130_fd_sc_hd__xor2_1
XFILLER_86_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2707 U$$4214/A1 U$$2707/A2 U$$3942/A1 U$$2707/B2 VGND VGND VPWR VPWR U$$2708/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2718 U$$2718/A U$$2734/B VGND VGND VPWR VPWR U$$2718/X sky130_fd_sc_hd__xor2_1
XFILLER_34_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2729 U$$2866/A1 U$$2729/A2 _612_/Q U$$2729/B2 VGND VGND VPWR VPWR U$$2730/A sky130_fd_sc_hd__a22o_1
XFILLER_160_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_413_ _541_/CLK _413_/D VGND VGND VPWR VPWR _413_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_775 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_344_ _475_/CLK _344_/D VGND VGND VPWR VPWR _344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_747 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_275_ _523_/CLK _275_/D VGND VGND VPWR VPWR _275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_482 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_80_0 dadda_fa_6_80_0/A dadda_fa_6_80_0/B dadda_fa_6_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_81_0/B dadda_fa_7_80_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_10_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_96_0 dadda_fa_3_96_0/A dadda_fa_3_96_0/B dadda_fa_3_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_0/B dadda_fa_4_96_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater906 U$$4382/B VGND VGND VPWR VPWR U$$4383/A sky130_fd_sc_hd__buf_6
XFILLER_111_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater917 U$$4247/A VGND VGND VPWR VPWR U$$4215/B sky130_fd_sc_hd__buf_8
Xrepeater928 _675_/Q VGND VGND VPWR VPWR U$$4070/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_58_5 dadda_fa_2_58_5/A dadda_fa_2_58_5/B dadda_fa_2_58_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_2/A dadda_fa_4_58_0/A sky130_fd_sc_hd__fa_2
Xrepeater939 U$$3764/B VGND VGND VPWR VPWR U$$3740/B sky130_fd_sc_hd__buf_6
XFILLER_209_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3920 _590_/Q U$$3932/A2 U$$4194/B1 U$$3932/B2 VGND VGND VPWR VPWR U$$3921/A sky130_fd_sc_hd__a22o_1
XFILLER_209_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3931 U$$3931/A U$$3935/B VGND VGND VPWR VPWR U$$3931/X sky130_fd_sc_hd__xor2_1
XU$$3942 U$$3942/A1 U$$3968/A2 U$$4218/A1 U$$3968/B2 VGND VGND VPWR VPWR U$$3943/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3953 U$$3953/A U$$3973/A VGND VGND VPWR VPWR U$$3953/X sky130_fd_sc_hd__xor2_1
XU$$3964 U$$4238/A1 U$$3970/A2 U$$4238/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3965/A
+ sky130_fd_sc_hd__a22o_1
XU$$3975 U$$4084/B VGND VGND VPWR VPWR U$$3975/Y sky130_fd_sc_hd__inv_1
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3986 U$$3986/A U$$3994/B VGND VGND VPWR VPWR U$$3986/X sky130_fd_sc_hd__xor2_1
XU$$3997 _560_/Q U$$4035/A2 U$$4273/A1 U$$4081/B2 VGND VGND VPWR VPWR U$$3998/A sky130_fd_sc_hd__a22o_1
XFILLER_127_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$180 U$$180/A U$$180/B VGND VGND VPWR VPWR U$$180/X sky130_fd_sc_hd__xor2_1
XU$$191 U$$54/A1 U$$219/A2 U$$56/A1 U$$219/B2 VGND VGND VPWR VPWR U$$192/A sky130_fd_sc_hd__a22o_1
XFILLER_205_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput266 _276_/Q VGND VGND VPWR VPWR o[108] sky130_fd_sc_hd__buf_2
Xrepeater1080 U$$1780/A VGND VGND VPWR VPWR U$$1773/B sky130_fd_sc_hd__buf_8
XFILLER_99_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput277 _286_/Q VGND VGND VPWR VPWR o[118] sky130_fd_sc_hd__buf_2
XFILLER_134_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1091 _639_/Q VGND VGND VPWR VPWR U$$1636/B sky130_fd_sc_hd__buf_6
XFILLER_114_563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput288 _180_/Q VGND VGND VPWR VPWR o[12] sky130_fd_sc_hd__buf_2
Xoutput299 _190_/Q VGND VGND VPWR VPWR o[22] sky130_fd_sc_hd__buf_2
XFILLER_99_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_60_5 U$$3984/X U$$4117/X U$$4141/B VGND VGND VPWR VPWR dadda_fa_2_61_2/A
+ dadda_fa_2_60_5/A sky130_fd_sc_hd__fa_1
XFILLER_101_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_53_4 U$$1975/X U$$2108/X U$$2241/X VGND VGND VPWR VPWR dadda_fa_2_54_1/CIN
+ dadda_fa_2_53_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_46_3 U$$1296/X U$$1429/X U$$1562/X VGND VGND VPWR VPWR dadda_fa_2_47_2/CIN
+ dadda_fa_2_46_5/A sky130_fd_sc_hd__fa_1
XFILLER_43_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_23_2 dadda_fa_4_23_2/A dadda_fa_4_23_2/B dadda_fa_4_23_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/CIN dadda_fa_5_23_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_16_1 U$$1103/X U$$1195/B input164/X VGND VGND VPWR VPWR dadda_fa_5_17_0/B
+ dadda_fa_5_16_1/B sky130_fd_sc_hd__fa_1
XFILLER_196_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_992 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_20 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3205 U$$4436/B1 U$$3285/A2 U$$4301/B1 U$$3285/B2 VGND VGND VPWR VPWR U$$3206/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_101_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3216 U$$3216/A U$$3218/B VGND VGND VPWR VPWR U$$3216/X sky130_fd_sc_hd__xor2_1
XFILLER_47_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3227 U$$3362/B1 U$$3231/A2 U$$3229/A1 U$$3231/B2 VGND VGND VPWR VPWR U$$3228/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3238 U$$3238/A U$$3286/B VGND VGND VPWR VPWR U$$3238/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2504 U$$2641/A1 U$$2550/A2 U$$2641/B1 U$$2550/B2 VGND VGND VPWR VPWR U$$2505/A
+ sky130_fd_sc_hd__a22o_1
XU$$3249 _597_/Q U$$3273/A2 _598_/Q U$$3273/B2 VGND VGND VPWR VPWR U$$3250/A sky130_fd_sc_hd__a22o_1
XU$$2515 U$$2515/A U$$2517/B VGND VGND VPWR VPWR U$$2515/X sky130_fd_sc_hd__xor2_1
XU$$2526 U$$334/A1 U$$2530/A2 U$$62/A1 U$$2530/B2 VGND VGND VPWR VPWR U$$2527/A sky130_fd_sc_hd__a22o_1
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2537 U$$2537/A U$$2567/B VGND VGND VPWR VPWR U$$2537/X sky130_fd_sc_hd__xor2_1
XU$$1803 U$$20/B1 U$$1843/A2 U$$2077/B1 U$$1843/B2 VGND VGND VPWR VPWR U$$1804/A sky130_fd_sc_hd__a22o_1
XU$$2548 U$$80/B1 U$$2550/A2 U$$906/A1 U$$2550/B2 VGND VGND VPWR VPWR U$$2549/A sky130_fd_sc_hd__a22o_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2559 U$$2559/A U$$2603/A VGND VGND VPWR VPWR U$$2559/X sky130_fd_sc_hd__xor2_1
XFILLER_62_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1814 U$$1814/A U$$1874/B VGND VGND VPWR VPWR U$$1814/X sky130_fd_sc_hd__xor2_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1825 U$$3056/B1 U$$1855/A2 U$$731/A1 U$$1855/B2 VGND VGND VPWR VPWR U$$1826/A
+ sky130_fd_sc_hd__a22o_1
XU$$1836 U$$1836/A U$$1844/B VGND VGND VPWR VPWR U$$1836/X sky130_fd_sc_hd__xor2_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1847 U$$3217/A1 U$$1915/A2 U$$4450/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1848/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1858 U$$1858/A U$$1870/B VGND VGND VPWR VPWR U$$1858/X sky130_fd_sc_hd__xor2_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1869 U$$2963/B1 U$$1785/X U$$90/A1 U$$1786/X VGND VGND VPWR VPWR U$$1870/A sky130_fd_sc_hd__a22o_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_79 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_327_ _455_/CLK _327_/D VGND VGND VPWR VPWR _327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_258_ _379_/CLK _258_/D VGND VGND VPWR VPWR _258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_189_ _189_/CLK _189_/D VGND VGND VPWR VPWR _189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_70_4 dadda_fa_2_70_4/A dadda_fa_2_70_4/B dadda_fa_2_70_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/CIN dadda_fa_3_70_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_97_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_63_3 dadda_fa_2_63_3/A dadda_fa_2_63_3/B dadda_fa_2_63_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/B dadda_fa_3_63_3/B sky130_fd_sc_hd__fa_1
Xrepeater703 U$$3932/B2 VGND VGND VPWR VPWR U$$3916/B2 sky130_fd_sc_hd__buf_4
Xrepeater714 U$$3805/B2 VGND VGND VPWR VPWR U$$3795/B2 sky130_fd_sc_hd__buf_4
XFILLER_42_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater725 U$$3567/X VGND VGND VPWR VPWR U$$3674/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_56_2 dadda_fa_2_56_2/A dadda_fa_2_56_2/B dadda_fa_2_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/A dadda_fa_3_56_3/A sky130_fd_sc_hd__fa_1
Xrepeater736 U$$3378/B2 VGND VGND VPWR VPWR U$$3320/B2 sky130_fd_sc_hd__clkbuf_8
Xrepeater747 U$$3273/B2 VGND VGND VPWR VPWR U$$3263/B2 sky130_fd_sc_hd__buf_4
Xrepeater758 U$$3019/X VGND VGND VPWR VPWR U$$3148/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_33_1 dadda_fa_5_33_1/A dadda_fa_5_33_1/B dadda_fa_5_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_34_0/B dadda_fa_7_33_0/A sky130_fd_sc_hd__fa_1
Xrepeater769 U$$398/B2 VGND VGND VPWR VPWR U$$334/B2 sky130_fd_sc_hd__buf_6
XU$$4440 U$$4440/A1 U$$4388/X U$$4442/A1 U$$4480/B2 VGND VGND VPWR VPWR U$$4441/A
+ sky130_fd_sc_hd__a22o_1
XU$$4451 U$$4451/A U$$4451/B VGND VGND VPWR VPWR U$$4451/X sky130_fd_sc_hd__xor2_1
XFILLER_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4462 U$$4462/A1 U$$4388/X U$$4464/A1 U$$4468/B2 VGND VGND VPWR VPWR U$$4463/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_1 dadda_fa_2_49_1/A dadda_fa_2_49_1/B dadda_fa_2_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_0/CIN dadda_fa_3_49_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_77_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4473 U$$4473/A U$$4473/B VGND VGND VPWR VPWR U$$4473/X sky130_fd_sc_hd__xor2_1
XU$$4484 U$$4484/A1 U$$4388/X U$$4486/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4485/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3750 U$$3750/A U$$3760/B VGND VGND VPWR VPWR U$$3750/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_26_0 dadda_fa_5_26_0/A dadda_fa_5_26_0/B dadda_fa_5_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_27_0/A dadda_fa_6_26_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_77_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4495 U$$4495/A U$$4495/B VGND VGND VPWR VPWR U$$4495/X sky130_fd_sc_hd__xor2_1
XU$$3761 U$$4444/B1 U$$3777/A2 U$$4448/A1 U$$3777/B2 VGND VGND VPWR VPWR U$$3762/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3772 U$$3772/A U$$3816/B VGND VGND VPWR VPWR U$$3772/X sky130_fd_sc_hd__xor2_1
XFILLER_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3783 U$$3783/A1 U$$3795/A2 U$$3783/B1 U$$3795/B2 VGND VGND VPWR VPWR U$$3784/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3794 U$$3794/A U$$3804/B VGND VGND VPWR VPWR U$$3794/X sky130_fd_sc_hd__xor2_1
XFILLER_52_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_100_0 dadda_fa_5_100_0/A dadda_fa_5_100_0/B dadda_fa_5_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_101_0/A dadda_fa_6_100_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_146_496 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_308 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_51_1 U$$508/X U$$641/X U$$774/X VGND VGND VPWR VPWR dadda_fa_2_52_0/CIN
+ dadda_fa_2_51_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_60_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$905 U$$905/A U$$907/B VGND VGND VPWR VPWR U$$905/X sky130_fd_sc_hd__xor2_1
XFILLER_21_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$916 U$$916/A1 U$$956/A2 U$$916/B1 U$$956/B2 VGND VGND VPWR VPWR U$$917/A sky130_fd_sc_hd__a22o_1
XFILLER_84_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$927 U$$927/A U$$935/B VGND VGND VPWR VPWR U$$927/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_44_0 U$$95/X U$$228/X U$$361/X VGND VGND VPWR VPWR dadda_fa_2_45_2/B dadda_fa_2_44_4/B
+ sky130_fd_sc_hd__fa_1
XFILLER_71_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$938 U$$938/A1 U$$826/X U$$938/B1 U$$827/X VGND VGND VPWR VPWR U$$939/A sky130_fd_sc_hd__a22o_1
XU$$949 U$$949/A U$$951/B VGND VGND VPWR VPWR U$$949/X sky130_fd_sc_hd__xor2_1
XFILLER_141_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_399 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_706 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_923 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_80_3 dadda_fa_3_80_3/A dadda_fa_3_80_3/B dadda_fa_3_80_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_1/B dadda_fa_4_80_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_999 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_73_2 dadda_fa_3_73_2/A dadda_fa_3_73_2/B dadda_fa_3_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_1/A dadda_fa_4_73_2/B sky130_fd_sc_hd__fa_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_66_1 dadda_fa_3_66_1/A dadda_fa_3_66_1/B dadda_fa_3_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_0/CIN dadda_fa_4_66_2/A sky130_fd_sc_hd__fa_1
XFILLER_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_43_0 dadda_fa_6_43_0/A dadda_fa_6_43_0/B dadda_fa_6_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_44_0/B dadda_fa_7_43_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_59_0 dadda_fa_3_59_0/A dadda_fa_3_59_0/B dadda_fa_3_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_0/B dadda_fa_4_59_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3002 U$$3002/A U$$3008/B VGND VGND VPWR VPWR U$$3002/X sky130_fd_sc_hd__xor2_1
XFILLER_207_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3013 U$$3014/A VGND VGND VPWR VPWR U$$3013/Y sky130_fd_sc_hd__inv_1
XFILLER_46_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3024 U$$556/B1 U$$3054/A2 U$$3024/B1 U$$3054/B2 VGND VGND VPWR VPWR U$$3025/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3035 U$$3035/A U$$3049/B VGND VGND VPWR VPWR U$$3035/X sky130_fd_sc_hd__xor2_1
XFILLER_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2301 U$$2301/A U$$2303/B VGND VGND VPWR VPWR U$$2301/X sky130_fd_sc_hd__xor2_1
XU$$3046 U$$3181/B1 U$$3046/A2 U$$3046/B1 U$$3046/B2 VGND VGND VPWR VPWR U$$3047/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3057 U$$3057/A U$$3065/B VGND VGND VPWR VPWR U$$3057/X sky130_fd_sc_hd__xor2_1
XU$$2312 U$$940/B1 U$$2318/A2 U$$3273/A1 U$$2318/B2 VGND VGND VPWR VPWR U$$2313/A
+ sky130_fd_sc_hd__a22o_1
XU$$2323 U$$2323/A U$$2328/A VGND VGND VPWR VPWR U$$2323/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_102_2 dadda_fa_4_102_2/A dadda_fa_4_102_2/B dadda_fa_4_102_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/CIN dadda_fa_5_102_1/CIN sky130_fd_sc_hd__fa_1
XU$$3068 U$$4436/B1 U$$3148/A2 U$$4301/B1 U$$3148/B2 VGND VGND VPWR VPWR U$$3069/A
+ sky130_fd_sc_hd__a22o_1
XU$$2334 U$$2332/B _649_/Q _650_/Q U$$2329/Y VGND VGND VPWR VPWR U$$2334/X sky130_fd_sc_hd__a22o_1
XFILLER_207_478 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1600 U$$1600/A U$$1642/B VGND VGND VPWR VPWR U$$1600/X sky130_fd_sc_hd__xor2_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3079 U$$3079/A U$$3083/B VGND VGND VPWR VPWR U$$3079/X sky130_fd_sc_hd__xor2_1
XU$$2345 U$$2345/A1 U$$2367/A2 U$$2895/A1 U$$2367/B2 VGND VGND VPWR VPWR U$$2346/A
+ sky130_fd_sc_hd__a22o_1
XU$$2356 U$$2356/A U$$2388/B VGND VGND VPWR VPWR U$$2356/X sky130_fd_sc_hd__xor2_1
XFILLER_90_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1611 U$$2431/B1 U$$1635/A2 U$$2435/A1 U$$1635/B2 VGND VGND VPWR VPWR U$$1612/A
+ sky130_fd_sc_hd__a22o_1
XU$$1622 U$$1622/A U$$1628/B VGND VGND VPWR VPWR U$$1622/X sky130_fd_sc_hd__xor2_1
XU$$2367 U$$2641/A1 U$$2367/A2 U$$2641/B1 U$$2367/B2 VGND VGND VPWR VPWR U$$2368/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2378 U$$2378/A U$$2418/B VGND VGND VPWR VPWR U$$2378/X sky130_fd_sc_hd__xor2_1
XFILLER_90_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1633 U$$946/B1 U$$1635/A2 U$$950/A1 U$$1635/B2 VGND VGND VPWR VPWR U$$1634/A sky130_fd_sc_hd__a22o_1
XU$$1644 _639_/Q VGND VGND VPWR VPWR U$$1644/Y sky130_fd_sc_hd__inv_1
XU$$2389 U$$334/A1 U$$2395/A2 U$$334/B1 U$$2395/B2 VGND VGND VPWR VPWR U$$2390/A sky130_fd_sc_hd__a22o_1
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1655 U$$1655/A U$$1687/B VGND VGND VPWR VPWR U$$1655/X sky130_fd_sc_hd__xor2_1
XFILLER_163_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1666 U$$20/B1 U$$1718/A2 U$$981/B1 U$$1718/B2 VGND VGND VPWR VPWR U$$1667/A sky130_fd_sc_hd__a22o_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1677 U$$1677/A U$$1719/B VGND VGND VPWR VPWR U$$1677/X sky130_fd_sc_hd__xor2_1
XFILLER_203_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$408_1761 VGND VGND VPWR VPWR U$$408_1761/HI U$$408/B1 sky130_fd_sc_hd__conb_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1688 U$$3056/B1 U$$1736/A2 U$$731/A1 U$$1736/B2 VGND VGND VPWR VPWR U$$1689/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1699 U$$1699/A U$$1719/B VGND VGND VPWR VPWR U$$1699/X sky130_fd_sc_hd__xor2_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_116_0 dadda_fa_7_116_0/A dadda_fa_7_116_0/B dadda_fa_7_116_0/CIN VGND
+ VGND VPWR VPWR _541_/D _412_/D sky130_fd_sc_hd__fa_1
XFILLER_204_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4457_1807 VGND VGND VPWR VPWR U$$4457_1807/HI U$$4457/B sky130_fd_sc_hd__conb_1
XFILLER_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_1125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1035 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_308 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_61_0 dadda_fa_2_61_0/A dadda_fa_2_61_0/B dadda_fa_2_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_0/B dadda_fa_3_61_2/B sky130_fd_sc_hd__fa_1
Xrepeater500 U$$3155/X VGND VGND VPWR VPWR U$$3273/A2 sky130_fd_sc_hd__clkbuf_8
Xfinal_adder.U$$307 final_adder.U$$306/A final_adder.U$$229/X final_adder.U$$231/X
+ VGND VGND VPWR VPWR final_adder.U$$307/X sky130_fd_sc_hd__a21o_1
Xrepeater511 U$$2973/A2 VGND VGND VPWR VPWR U$$2929/A2 sky130_fd_sc_hd__buf_4
XFILLER_97_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater522 U$$408/A2 VGND VGND VPWR VPWR U$$398/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$329 final_adder.U$$328/A final_adder.U$$273/X final_adder.U$$275/X
+ VGND VGND VPWR VPWR final_adder.U$$329/X sky130_fd_sc_hd__a21o_1
XFILLER_69_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater533 U$$2874/A2 VGND VGND VPWR VPWR U$$2866/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater544 U$$2470/X VGND VGND VPWR VPWR U$$2566/A2 sky130_fd_sc_hd__buf_6
Xrepeater555 U$$2463/A2 VGND VGND VPWR VPWR U$$2423/A2 sky130_fd_sc_hd__buf_4
Xrepeater566 U$$2196/X VGND VGND VPWR VPWR U$$2318/A2 sky130_fd_sc_hd__buf_4
XFILLER_211_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater577 U$$2010/A2 VGND VGND VPWR VPWR U$$1982/A2 sky130_fd_sc_hd__buf_6
Xrepeater588 U$$1909/A2 VGND VGND VPWR VPWR U$$1915/A2 sky130_fd_sc_hd__buf_6
XU$$4270 U$$4270/A U$$4298/B VGND VGND VPWR VPWR U$$4270/X sky130_fd_sc_hd__xor2_1
XU$$4281 U$$4418/A1 U$$4327/A2 U$$4418/B1 U$$4319/B2 VGND VGND VPWR VPWR U$$4282/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater599 U$$1553/A2 VGND VGND VPWR VPWR U$$1557/A2 sky130_fd_sc_hd__buf_6
XU$$4292 U$$4292/A U$$4296/B VGND VGND VPWR VPWR U$$4292/X sky130_fd_sc_hd__xor2_1
XFILLER_93_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3580 _557_/Q U$$3628/A2 U$$4404/A1 U$$3628/B2 VGND VGND VPWR VPWR U$$3581/A sky130_fd_sc_hd__a22o_1
XU$$3591 U$$3591/A U$$3637/B VGND VGND VPWR VPWR U$$3591/X sky130_fd_sc_hd__xor2_1
XFILLER_179_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2890 U$$2890/A U$$2928/B VGND VGND VPWR VPWR U$$2890/X sky130_fd_sc_hd__xor2_1
XFILLER_178_330 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_90_2 dadda_fa_4_90_2/A dadda_fa_4_90_2/B dadda_fa_4_90_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/CIN dadda_fa_5_90_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_83_1 dadda_fa_4_83_1/A dadda_fa_4_83_1/B dadda_fa_4_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/B dadda_fa_5_83_1/B sky130_fd_sc_hd__fa_1
XFILLER_134_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_60_0 dadda_fa_7_60_0/A dadda_fa_7_60_0/B dadda_fa_7_60_0/CIN VGND VGND
+ VPWR VPWR _485_/D _356_/D sky130_fd_sc_hd__fa_1
XFILLER_135_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_76_0 dadda_fa_4_76_0/A dadda_fa_4_76_0/B dadda_fa_4_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/A dadda_fa_5_76_1/A sky130_fd_sc_hd__fa_1
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_661_ _674_/CLK _661_/D VGND VGND VPWR VPWR _661_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$702 U$$702/A U$$726/B VGND VGND VPWR VPWR U$$702/X sky130_fd_sc_hd__xor2_1
XU$$713 U$$848/B1 U$$765/A2 U$$715/A1 U$$765/B2 VGND VGND VPWR VPWR U$$714/A sky130_fd_sc_hd__a22o_1
XFILLER_44_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$724 U$$724/A U$$726/B VGND VGND VPWR VPWR U$$724/X sky130_fd_sc_hd__xor2_1
XFILLER_90_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_592_ _596_/CLK _592_/D VGND VGND VPWR VPWR _592_/Q sky130_fd_sc_hd__dfxtp_1
XU$$735 U$$48/B1 U$$747/A2 U$$874/A1 U$$747/B2 VGND VGND VPWR VPWR U$$736/A sky130_fd_sc_hd__a22o_1
XFILLER_72_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$746 U$$746/A U$$748/B VGND VGND VPWR VPWR U$$746/X sky130_fd_sc_hd__xor2_1
XFILLER_56_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$757 U$$757/A1 U$$795/A2 U$$759/A1 U$$795/B2 VGND VGND VPWR VPWR U$$758/A sky130_fd_sc_hd__a22o_1
XFILLER_43_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$768 U$$768/A U$$816/B VGND VGND VPWR VPWR U$$768/X sky130_fd_sc_hd__xor2_1
XU$$779 U$$914/B1 U$$783/A2 U$$916/B1 U$$783/B2 VGND VGND VPWR VPWR U$$780/A sky130_fd_sc_hd__a22o_1
XFILLER_147_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1602 _565_/Q VGND VGND VPWR VPWR U$$3046/B1 sky130_fd_sc_hd__buf_8
XANTENNA_7 _472_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1613 U$$2494/B1 VGND VGND VPWR VPWR U$$30/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1624 U$$4273/B1 VGND VGND VPWR VPWR U$$3453/A1 sky130_fd_sc_hd__buf_6
Xrepeater1635 _561_/Q VGND VGND VPWR VPWR U$$4410/A1 sky130_fd_sc_hd__buf_4
Xrepeater1646 U$$22/A1 VGND VGND VPWR VPWR U$$707/A1 sky130_fd_sc_hd__clkbuf_4
Xrepeater1657 U$$840/B1 VGND VGND VPWR VPWR U$$705/A1 sky130_fd_sc_hd__buf_6
Xrepeater1668 _557_/Q VGND VGND VPWR VPWR U$$4402/A1 sky130_fd_sc_hd__buf_4
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1679 U$$2343/A1 VGND VGND VPWR VPWR U$$14/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_40_5 dadda_fa_2_40_5/A dadda_fa_2_40_5/B dadda_fa_2_40_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_41_2/A dadda_fa_4_40_0/A sky130_fd_sc_hd__fa_2
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_33_4 U$$1669/X U$$1802/X U$$1935/X VGND VGND VPWR VPWR dadda_fa_3_34_1/CIN
+ dadda_fa_3_33_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2120 U$$2120/A U$$2144/B VGND VGND VPWR VPWR U$$2120/X sky130_fd_sc_hd__xor2_1
XU$$2131 U$$3638/A1 U$$2135/A2 U$$3503/A1 U$$2135/B2 VGND VGND VPWR VPWR U$$2132/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2142 U$$2142/A U$$2174/B VGND VGND VPWR VPWR U$$2142/X sky130_fd_sc_hd__xor2_1
XU$$2153 U$$3521/B1 U$$2189/A2 U$$3386/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2154/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2164 U$$2164/A U$$2186/B VGND VGND VPWR VPWR U$$2164/X sky130_fd_sc_hd__xor2_1
XU$$2175 U$$940/B1 U$$2185/A2 U$$3273/A1 U$$2185/B2 VGND VGND VPWR VPWR U$$2176/A
+ sky130_fd_sc_hd__a22o_1
XU$$1430 U$$882/A1 U$$1478/A2 U$$3213/A1 U$$1478/B2 VGND VGND VPWR VPWR U$$1431/A
+ sky130_fd_sc_hd__a22o_1
XU$$1441 U$$1441/A U$$1443/B VGND VGND VPWR VPWR U$$1441/X sky130_fd_sc_hd__xor2_1
XU$$2186 U$$2186/A U$$2186/B VGND VGND VPWR VPWR U$$2186/X sky130_fd_sc_hd__xor2_1
XFILLER_179_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2197 U$$2195/B _647_/Q _648_/Q U$$2192/Y VGND VGND VPWR VPWR U$$2197/X sky130_fd_sc_hd__a22o_1
XU$$1452 U$$82/A1 U$$1478/A2 U$$3096/B1 U$$1478/B2 VGND VGND VPWR VPWR U$$1453/A sky130_fd_sc_hd__a22o_1
XU$$1463 U$$1463/A U$$1475/B VGND VGND VPWR VPWR U$$1463/X sky130_fd_sc_hd__xor2_1
XFILLER_15_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1474 U$$924/B1 U$$1474/A2 U$$2435/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1475/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1485 U$$1485/A U$$1487/B VGND VGND VPWR VPWR U$$1485/X sky130_fd_sc_hd__xor2_1
XU$$1496 U$$948/A1 U$$1500/A2 U$$948/B1 U$$1500/B2 VGND VGND VPWR VPWR U$$1497/A sky130_fd_sc_hd__a22o_1
XFILLER_163_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_93_0 dadda_fa_5_93_0/A dadda_fa_5_93_0/B dadda_fa_5_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_94_0/A dadda_fa_6_93_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_78_6 U$$3621/X U$$3754/X U$$3887/X VGND VGND VPWR VPWR dadda_fa_2_79_2/B
+ dadda_fa_2_78_5/B sky130_fd_sc_hd__fa_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4511_1834 VGND VGND VPWR VPWR U$$4511_1834/HI U$$4511/B sky130_fd_sc_hd__conb_1
XFILLER_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1095 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$104 _528_/Q _400_/Q VGND VGND VPWR VPWR final_adder.U$$599/B1 final_adder.U$$726/A
+ sky130_fd_sc_hd__ha_2
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$115 _539_/Q _411_/Q VGND VGND VPWR VPWR final_adder.U$$243/B1 final_adder.U$$737/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$126 _550_/Q _422_/Q VGND VGND VPWR VPWR final_adder.U$$621/B1 final_adder.U$$748/A
+ sky130_fd_sc_hd__ha_2
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$137 final_adder.U$$9/SUM final_adder.U$$8/COUT final_adder.U$$9/COUT
+ VGND VGND VPWR VPWR final_adder.U$$137/X sky130_fd_sc_hd__a21o_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$148 final_adder.U$$643/A final_adder.U$$642/A VGND VGND VPWR VPWR
+ final_adder.U$$266/B sky130_fd_sc_hd__and2_1
XFILLER_211_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$159 final_adder.U$$653/A final_adder.U$$525/B1 final_adder.U$$159/B1
+ VGND VGND VPWR VPWR final_adder.U$$159/X sky130_fd_sc_hd__a21o_1
XFILLER_73_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater385 U$$1065/A2 VGND VGND VPWR VPWR U$$995/A2 sky130_fd_sc_hd__buf_4
XFILLER_54_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater396 U$$896/A2 VGND VGND VPWR VPWR U$$906/A2 sky130_fd_sc_hd__buf_4
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_420 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_102_1 U$$4467/X input132/X dadda_fa_3_102_1/CIN VGND VGND VPWR VPWR dadda_fa_4_103_0/CIN
+ dadda_fa_4_102_2/A sky130_fd_sc_hd__fa_1
XFILLER_190_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_959 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput100 b[41] VGND VGND VPWR VPWR _593_/D sky130_fd_sc_hd__clkbuf_1
Xinput111 b[51] VGND VGND VPWR VPWR _603_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput122 b[61] VGND VGND VPWR VPWR _613_/D sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_6_123_0 dadda_fa_6_123_0/A dadda_fa_6_123_0/B dadda_fa_6_123_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_124_0/B dadda_fa_7_123_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput133 c[103] VGND VGND VPWR VPWR input133/X sky130_fd_sc_hd__buf_2
XFILLER_62_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput144 c[113] VGND VGND VPWR VPWR input144/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_66_4 U$$1735/X U$$1868/X U$$2001/X VGND VGND VPWR VPWR dadda_fa_1_67_6/CIN
+ dadda_fa_1_66_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput155 c[123] VGND VGND VPWR VPWR input155/X sky130_fd_sc_hd__clkbuf_1
XTAP_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 c[18] VGND VGND VPWR VPWR input166/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput177 c[28] VGND VGND VPWR VPWR input177/X sky130_fd_sc_hd__clkbuf_1
XTAP_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_43_3 dadda_fa_3_43_3/A dadda_fa_3_43_3/B dadda_fa_3_43_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_1/B dadda_fa_4_43_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 c[38] VGND VGND VPWR VPWR input188/X sky130_fd_sc_hd__clkbuf_4
XTAP_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput199 c[48] VGND VGND VPWR VPWR input199/X sky130_fd_sc_hd__buf_2
XFILLER_76_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$660 final_adder.U$$660/A final_adder.U$$660/B VGND VGND VPWR VPWR
+ _206_/D sky130_fd_sc_hd__xor2_1
XTAP_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$671 final_adder.U$$671/A final_adder.U$$671/B VGND VGND VPWR VPWR
+ _217_/D sky130_fd_sc_hd__xor2_1
XTAP_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$510 U$$510/A U$$518/B VGND VGND VPWR VPWR U$$510/X sky130_fd_sc_hd__xor2_1
X_644_ _648_/CLK _644_/D VGND VGND VPWR VPWR _644_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$682 final_adder.U$$682/A final_adder.U$$682/B VGND VGND VPWR VPWR
+ _228_/D sky130_fd_sc_hd__xor2_1
XTAP_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_36_2 dadda_fa_3_36_2/A dadda_fa_3_36_2/B dadda_fa_3_36_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_1/A dadda_fa_4_36_2/B sky130_fd_sc_hd__fa_1
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$521 U$$658/A1 U$$545/A2 U$$658/B1 U$$545/B2 VGND VGND VPWR VPWR U$$522/A sky130_fd_sc_hd__a22o_1
XFILLER_205_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$532 U$$532/A U$$532/B VGND VGND VPWR VPWR U$$532/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$693 final_adder.U$$693/A final_adder.U$$693/B VGND VGND VPWR VPWR
+ _239_/D sky130_fd_sc_hd__xor2_4
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$543 U$$678/B1 U$$545/A2 U$$545/A1 U$$545/B2 VGND VGND VPWR VPWR U$$544/A sky130_fd_sc_hd__a22o_1
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_29_1 U$$1927/X input178/X dadda_fa_3_29_1/CIN VGND VGND VPWR VPWR dadda_fa_4_30_0/CIN
+ dadda_fa_4_29_2/A sky130_fd_sc_hd__fa_1
XU$$554 U$$554/A1 U$$600/A2 U$$828/B1 U$$600/B2 VGND VGND VPWR VPWR U$$555/A sky130_fd_sc_hd__a22o_1
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_575_ _575_/CLK _575_/D VGND VGND VPWR VPWR _575_/Q sky130_fd_sc_hd__dfxtp_4
XU$$565 U$$565/A U$$589/B VGND VGND VPWR VPWR U$$565/X sky130_fd_sc_hd__xor2_1
XFILLER_60_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$576 U$$848/B1 U$$600/A2 U$$715/A1 U$$600/B2 VGND VGND VPWR VPWR U$$577/A sky130_fd_sc_hd__a22o_1
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$587 U$$587/A U$$627/B VGND VGND VPWR VPWR U$$587/X sky130_fd_sc_hd__xor2_1
XU$$598 U$$733/B1 U$$600/A2 U$$600/A1 U$$600/B2 VGND VGND VPWR VPWR U$$599/A sky130_fd_sc_hd__a22o_1
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1410 _589_/Q VGND VGND VPWR VPWR U$$4466/A1 sky130_fd_sc_hd__buf_2
Xrepeater1421 U$$3229/A1 VGND VGND VPWR VPWR U$$900/A1 sky130_fd_sc_hd__buf_6
XFILLER_160_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1432 U$$4323/A1 VGND VGND VPWR VPWR U$$3638/A1 sky130_fd_sc_hd__buf_6
XFILLER_158_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1443 U$$894/A1 VGND VGND VPWR VPWR U$$72/A1 sky130_fd_sc_hd__buf_6
Xrepeater1454 _583_/Q VGND VGND VPWR VPWR U$$3358/A1 sky130_fd_sc_hd__buf_6
XFILLER_119_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_88_5 dadda_fa_2_88_5/A dadda_fa_2_88_5/B dadda_fa_2_88_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_2/A dadda_fa_4_88_0/A sky130_fd_sc_hd__fa_2
Xrepeater1465 U$$4176/B1 VGND VGND VPWR VPWR U$$3902/B1 sky130_fd_sc_hd__buf_6
XFILLER_114_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1476 U$$749/A1 VGND VGND VPWR VPWR U$$747/B1 sky130_fd_sc_hd__buf_4
XFILLER_125_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1487 U$$3896/B1 VGND VGND VPWR VPWR U$$3213/A1 sky130_fd_sc_hd__buf_6
XFILLER_113_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1498 U$$4444/A1 VGND VGND VPWR VPWR U$$4168/B1 sky130_fd_sc_hd__buf_6
XFILLER_154_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_31_1 U$$468/X U$$601/X U$$734/X VGND VGND VPWR VPWR dadda_fa_3_32_1/A
+ dadda_fa_3_31_3/A sky130_fd_sc_hd__fa_1
XFILLER_39_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_24_0 U$$55/X U$$188/X U$$321/X VGND VGND VPWR VPWR dadda_fa_3_25_3/A dadda_fa_3_24_3/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1260 U$$1260/A U$$1288/B VGND VGND VPWR VPWR U$$1260/X sky130_fd_sc_hd__xor2_1
XU$$1271 U$$2641/A1 U$$1279/A2 U$$2641/B1 U$$1279/B2 VGND VGND VPWR VPWR U$$1272/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1282 U$$1282/A U$$1296/B VGND VGND VPWR VPWR U$$1282/X sky130_fd_sc_hd__xor2_1
XFILLER_206_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1293 U$$334/A1 U$$1323/A2 U$$334/B1 U$$1323/B2 VGND VGND VPWR VPWR U$$1294/A sky130_fd_sc_hd__a22o_1
XFILLER_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_118_1 dadda_fa_5_118_1/A dadda_fa_5_118_1/B dadda_ha_4_118_2/SUM VGND
+ VGND VPWR VPWR dadda_fa_6_119_0/B dadda_fa_7_118_0/A sky130_fd_sc_hd__fa_1
Xdadda_ha_1_84_6 U$$3766/X U$$3899/X VGND VGND VPWR VPWR dadda_fa_2_85_4/A dadda_fa_3_84_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_164_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_4 U$$2966/X U$$3099/X U$$3232/X VGND VGND VPWR VPWR dadda_fa_2_84_3/A
+ dadda_fa_2_83_5/B sky130_fd_sc_hd__fa_1
XFILLER_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_76_3 U$$2686/X U$$2819/X U$$2952/X VGND VGND VPWR VPWR dadda_fa_2_77_1/B
+ dadda_fa_2_76_4/B sky130_fd_sc_hd__fa_1
Xdadda_fa_4_53_2 dadda_fa_4_53_2/A dadda_fa_4_53_2/B dadda_fa_4_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/CIN dadda_fa_5_53_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_2 U$$3204/X U$$3337/X U$$3470/X VGND VGND VPWR VPWR dadda_fa_2_70_1/A
+ dadda_fa_2_69_4/A sky130_fd_sc_hd__fa_1
XFILLER_133_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_46_1 dadda_fa_4_46_1/A dadda_fa_4_46_1/B dadda_fa_4_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/B dadda_fa_5_46_1/B sky130_fd_sc_hd__fa_1
XFILLER_133_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_23_0 dadda_fa_7_23_0/A dadda_fa_7_23_0/B dadda_fa_7_23_0/CIN VGND VGND
+ VPWR VPWR _448_/D _319_/D sky130_fd_sc_hd__fa_1
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_39_0 dadda_fa_4_39_0/A dadda_fa_4_39_0/B dadda_fa_4_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/A dadda_fa_5_39_1/A sky130_fd_sc_hd__fa_1
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_216 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_227 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_238 _190_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_249 _195_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_360_ _491_/CLK _360_/D VGND VGND VPWR VPWR _360_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_291_ _615_/CLK _291_/D VGND VGND VPWR VPWR _291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_984 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_86_0_1857 VGND VGND VPWR VPWR dadda_fa_1_86_0/A dadda_fa_1_86_0_1857/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_123_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_71_2 U$$1346/X U$$1479/X U$$1612/X VGND VGND VPWR VPWR dadda_fa_1_72_7/B
+ dadda_fa_1_71_8/CIN sky130_fd_sc_hd__fa_1
XTAP_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_64_1 U$$534/X U$$667/X U$$800/X VGND VGND VPWR VPWR dadda_fa_1_65_5/CIN
+ dadda_fa_1_64_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_41_0 dadda_fa_3_41_0/A dadda_fa_3_41_0/B dadda_fa_3_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_0/B dadda_fa_4_41_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_92_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_57_0 U$$121/X U$$254/X U$$387/X VGND VGND VPWR VPWR dadda_fa_1_58_7/A
+ dadda_fa_1_57_8/B sky130_fd_sc_hd__fa_1
XTAP_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$340 U$$614/A1 U$$350/A2 U$$614/B1 U$$350/B2 VGND VGND VPWR VPWR U$$341/A sky130_fd_sc_hd__a22o_1
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_627_ _627_/CLK _627_/D VGND VGND VPWR VPWR _627_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$351 U$$351/A U$$351/B VGND VGND VPWR VPWR U$$351/X sky130_fd_sc_hd__xor2_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$362 U$$634/B1 U$$408/A2 U$$501/A1 U$$408/B2 VGND VGND VPWR VPWR U$$363/A sky130_fd_sc_hd__a22o_1
XFILLER_32_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$373 U$$373/A U$$383/B VGND VGND VPWR VPWR U$$373/X sky130_fd_sc_hd__xor2_1
XU$$384 U$$658/A1 U$$384/A2 U$$384/B1 U$$384/B2 VGND VGND VPWR VPWR U$$385/A sky130_fd_sc_hd__a22o_1
XU$$395 U$$395/A U$$410/A VGND VGND VPWR VPWR U$$395/X sky130_fd_sc_hd__xor2_1
X_558_ _558_/CLK _558_/D VGND VGND VPWR VPWR _558_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_489_ _491_/CLK _489_/D VGND VGND VPWR VPWR _489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_93_3 U$$4050/X U$$4183/X U$$4316/X VGND VGND VPWR VPWR dadda_fa_3_94_1/B
+ dadda_fa_3_93_3/B sky130_fd_sc_hd__fa_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1240 U$$944/A1 VGND VGND VPWR VPWR U$$942/B1 sky130_fd_sc_hd__buf_6
Xrepeater1251 U$$4504/A1 VGND VGND VPWR VPWR U$$4228/B1 sky130_fd_sc_hd__buf_6
Xrepeater1262 U$$3132/A1 VGND VGND VPWR VPWR U$$3952/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_86_2 input241/X dadda_fa_2_86_2/B dadda_fa_2_86_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_87_1/A dadda_fa_3_86_3/A sky130_fd_sc_hd__fa_1
Xrepeater1273 U$$2991/A1 VGND VGND VPWR VPWR U$$251/A1 sky130_fd_sc_hd__buf_8
XFILLER_99_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1284 U$$2715/A1 VGND VGND VPWR VPWR U$$658/B1 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_5_63_1 dadda_fa_5_63_1/A dadda_fa_5_63_1/B dadda_fa_5_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_64_0/B dadda_fa_7_63_0/A sky130_fd_sc_hd__fa_1
Xrepeater1295 U$$4355/B1 VGND VGND VPWR VPWR U$$4357/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_79_1 dadda_fa_2_79_1/A dadda_fa_2_79_1/B dadda_fa_2_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_0/CIN dadda_fa_3_79_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_56_0 dadda_fa_5_56_0/A dadda_fa_5_56_0/B dadda_fa_5_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_57_0/A dadda_fa_6_56_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_45_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_55_8 dadda_fa_1_55_8/A dadda_fa_1_55_8/B dadda_fa_1_55_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_56_3/A dadda_fa_3_55_0/A sky130_fd_sc_hd__fa_2
XFILLER_83_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_102_0 dadda_fa_2_102_0/A U$$2738/X U$$2871/X VGND VGND VPWR VPWR dadda_fa_3_103_2/A
+ dadda_fa_3_102_3/A sky130_fd_sc_hd__fa_1
XFILLER_208_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1090 U$$1090/A U$$1090/B VGND VGND VPWR VPWR U$$1090/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_74_0_1852 VGND VGND VPWR VPWR dadda_fa_0_74_0/A dadda_fa_0_74_0_1852/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_81_1 U$$1632/X U$$1765/X U$$1898/X VGND VGND VPWR VPWR dadda_fa_2_82_1/B
+ dadda_fa_2_81_4/A sky130_fd_sc_hd__fa_1
XFILLER_176_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_74_0 U$$1751/X U$$1884/X U$$2017/X VGND VGND VPWR VPWR dadda_fa_2_75_0/B
+ dadda_fa_2_74_3/B sky130_fd_sc_hd__fa_1
XFILLER_104_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3409 U$$3409/A U$$3425/A VGND VGND VPWR VPWR U$$3409/X sky130_fd_sc_hd__xor2_1
XFILLER_73_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2708 U$$2708/A U$$2708/B VGND VGND VPWR VPWR U$$2708/X sky130_fd_sc_hd__xor2_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2719 U$$2991/B1 U$$2729/A2 U$$2858/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2720/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_412_ _541_/CLK _412_/D VGND VGND VPWR VPWR _412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_343_ _343_/CLK _343_/D VGND VGND VPWR VPWR _343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_274_ _521_/CLK _274_/D VGND VGND VPWR VPWR _274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_96_1 dadda_fa_3_96_1/A dadda_fa_3_96_1/B dadda_fa_3_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_0/CIN dadda_fa_4_96_2/A sky130_fd_sc_hd__fa_1
XFILLER_182_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_73_0 dadda_fa_6_73_0/A dadda_fa_6_73_0/B dadda_fa_6_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_74_0/B dadda_fa_7_73_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_142_328 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_89_0 dadda_fa_3_89_0/A dadda_fa_3_89_0/B dadda_fa_3_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_0/B dadda_fa_4_89_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater907 U$$4350/B VGND VGND VPWR VPWR U$$4382/B sky130_fd_sc_hd__clkbuf_8
XFILLER_96_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater918 U$$4247/A VGND VGND VPWR VPWR U$$4175/B sky130_fd_sc_hd__buf_6
XFILLER_204_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater929 _675_/Q VGND VGND VPWR VPWR U$$4072/B sky130_fd_sc_hd__buf_6
XFILLER_110_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3910 U$$4456/B1 U$$3910/A2 U$$4323/A1 U$$3910/B2 VGND VGND VPWR VPWR U$$3911/A
+ sky130_fd_sc_hd__a22o_1
XU$$3921 U$$3921/A U$$3935/B VGND VGND VPWR VPWR U$$3921/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_118_0 dadda_fa_4_118_0/A U$$3834/X U$$3967/X VGND VGND VPWR VPWR dadda_fa_5_119_0/B
+ dadda_fa_5_118_1/A sky130_fd_sc_hd__fa_1
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3932 U$$3932/A1 U$$3932/A2 U$$918/B1 U$$3932/B2 VGND VGND VPWR VPWR U$$3933/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3943 U$$3943/A U$$3943/B VGND VGND VPWR VPWR U$$3943/X sky130_fd_sc_hd__xor2_1
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3954 U$$4502/A1 U$$3968/A2 U$$4504/A1 U$$3968/B2 VGND VGND VPWR VPWR U$$3955/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_5_5_0 U$$17/X U$$150/X VGND VGND VPWR VPWR dadda_fa_6_6_0/B dadda_fa_7_5_0/A
+ sky130_fd_sc_hd__ha_1
XU$$3965 U$$3965/A U$$3965/B VGND VGND VPWR VPWR U$$3965/X sky130_fd_sc_hd__xor2_1
XU$$3976 U$$4072/B U$$3976/B VGND VGND VPWR VPWR U$$3976/X sky130_fd_sc_hd__and2_1
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3987 U$$4259/B1 U$$4005/A2 U$$4400/A1 U$$4005/B2 VGND VGND VPWR VPWR U$$3988/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3998 U$$3998/A U$$4096/B VGND VGND VPWR VPWR U$$3998/X sky130_fd_sc_hd__xor2_1
XU$$170 U$$170/A U$$196/B VGND VGND VPWR VPWR U$$170/X sky130_fd_sc_hd__xor2_1
XU$$181 U$$44/A1 U$$181/A2 U$$46/A1 U$$181/B2 VGND VGND VPWR VPWR U$$182/A sky130_fd_sc_hd__a22o_1
XFILLER_127_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$192 U$$192/A U$$226/B VGND VGND VPWR VPWR U$$192/X sky130_fd_sc_hd__xor2_1
XFILLER_32_220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_448 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_91_0 U$$3115/X U$$3248/X U$$3381/X VGND VGND VPWR VPWR dadda_fa_3_92_0/B
+ dadda_fa_3_91_2/B sky130_fd_sc_hd__fa_1
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1070 U$$1918/A VGND VGND VPWR VPWR U$$1874/B sky130_fd_sc_hd__buf_8
Xoutput267 _277_/Q VGND VGND VPWR VPWR o[109] sky130_fd_sc_hd__buf_2
Xrepeater1081 U$$1780/A VGND VGND VPWR VPWR U$$1747/B sky130_fd_sc_hd__buf_8
Xrepeater1092 U$$1459/B VGND VGND VPWR VPWR U$$1425/B sky130_fd_sc_hd__buf_6
Xoutput278 _287_/Q VGND VGND VPWR VPWR o[119] sky130_fd_sc_hd__buf_2
Xoutput289 _181_/Q VGND VGND VPWR VPWR o[13] sky130_fd_sc_hd__buf_2
XFILLER_134_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_47_6 U$$2495/X U$$2628/X VGND VGND VPWR VPWR dadda_fa_2_48_3/B dadda_fa_3_47_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_101_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_60_6 input213/X dadda_fa_1_60_6/B dadda_fa_1_60_6/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_61_2/B dadda_fa_2_60_5/B sky130_fd_sc_hd__fa_1
XFILLER_114_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_53_5 U$$2374/X U$$2507/X U$$2640/X VGND VGND VPWR VPWR dadda_fa_2_54_2/A
+ dadda_fa_2_53_5/A sky130_fd_sc_hd__fa_1
XFILLER_114_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_46_4 U$$1695/X U$$1828/X U$$1961/X VGND VGND VPWR VPWR dadda_fa_2_47_3/A
+ dadda_fa_2_46_5/B sky130_fd_sc_hd__fa_1
XFILLER_15_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_16_2 dadda_fa_4_16_2/A dadda_fa_4_16_2/B dadda_ha_3_16_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_17_0/CIN dadda_fa_5_16_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_90_0 dadda_fa_7_90_0/A dadda_fa_7_90_0/B dadda_fa_7_90_0/CIN VGND VGND
+ VPWR VPWR _515_/D _386_/D sky130_fd_sc_hd__fa_1
XFILLER_177_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3206 U$$3206/A U$$3286/B VGND VGND VPWR VPWR U$$3206/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3217 U$$3217/A1 U$$3231/A2 U$$3354/B1 U$$3231/B2 VGND VGND VPWR VPWR U$$3218/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_1134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3228 U$$3228/A U$$3232/B VGND VGND VPWR VPWR U$$3228/X sky130_fd_sc_hd__xor2_1
XFILLER_47_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3239 U$$4472/A1 U$$3285/A2 U$$4474/A1 U$$3285/B2 VGND VGND VPWR VPWR U$$3240/A
+ sky130_fd_sc_hd__a22o_1
XU$$2505 U$$2505/A U$$2551/B VGND VGND VPWR VPWR U$$2505/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2516 U$$3475/A1 U$$2516/A2 U$$3475/B1 U$$2516/B2 VGND VGND VPWR VPWR U$$2517/A
+ sky130_fd_sc_hd__a22o_1
XU$$2527 U$$2527/A U$$2531/B VGND VGND VPWR VPWR U$$2527/X sky130_fd_sc_hd__xor2_1
XFILLER_64_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2538 U$$3769/B1 U$$2470/X U$$3771/B1 U$$2471/X VGND VGND VPWR VPWR U$$2539/A sky130_fd_sc_hd__a22o_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1804 U$$1804/A U$$1844/B VGND VGND VPWR VPWR U$$1804/X sky130_fd_sc_hd__xor2_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2549 U$$2549/A U$$2551/B VGND VGND VPWR VPWR U$$2549/X sky130_fd_sc_hd__xor2_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1815 U$$3320/B1 U$$1855/A2 U$$719/B1 U$$1855/B2 VGND VGND VPWR VPWR U$$1816/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1826 U$$1826/A U$$1874/B VGND VGND VPWR VPWR U$$1826/X sky130_fd_sc_hd__xor2_1
XU$$1837 U$$3618/A1 U$$1843/A2 U$$1976/A1 U$$1843/B2 VGND VGND VPWR VPWR U$$1838/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1848 U$$1848/A U$$1884/B VGND VGND VPWR VPWR U$$1848/X sky130_fd_sc_hd__xor2_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1859 U$$624/B1 U$$1859/A2 U$$491/A1 U$$1859/B2 VGND VGND VPWR VPWR U$$1860/A sky130_fd_sc_hd__a22o_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_326_ _454_/CLK _326_/D VGND VGND VPWR VPWR _326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_257_ _379_/CLK _257_/D VGND VGND VPWR VPWR _257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_188_ _207_/CLK _188_/D VGND VGND VPWR VPWR _188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_70_5 dadda_fa_2_70_5/A dadda_fa_2_70_5/B dadda_fa_2_70_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_2/A dadda_fa_4_70_0/A sky130_fd_sc_hd__fa_1
XFILLER_69_415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_63_4 dadda_fa_2_63_4/A dadda_fa_2_63_4/B dadda_fa_2_63_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/CIN dadda_fa_3_63_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater704 U$$3841/X VGND VGND VPWR VPWR U$$3932/B2 sky130_fd_sc_hd__buf_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater715 U$$3805/B2 VGND VGND VPWR VPWR U$$3777/B2 sky130_fd_sc_hd__buf_6
XFILLER_56_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater726 U$$3497/B2 VGND VGND VPWR VPWR U$$3479/B2 sky130_fd_sc_hd__buf_8
Xdadda_fa_2_56_3 dadda_fa_2_56_3/A dadda_fa_2_56_3/B dadda_fa_2_56_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/B dadda_fa_3_56_3/B sky130_fd_sc_hd__fa_1
Xrepeater737 U$$3378/B2 VGND VGND VPWR VPWR U$$3356/B2 sky130_fd_sc_hd__clkbuf_8
Xrepeater748 U$$3156/X VGND VGND VPWR VPWR U$$3273/B2 sky130_fd_sc_hd__clkbuf_8
XU$$4430 U$$4430/A1 U$$4388/X U$$4432/A1 U$$4430/B2 VGND VGND VPWR VPWR U$$4431/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater759 U$$2973/B2 VGND VGND VPWR VPWR U$$2929/B2 sky130_fd_sc_hd__buf_4
XU$$4441 U$$4441/A U$$4441/B VGND VGND VPWR VPWR U$$4441/X sky130_fd_sc_hd__xor2_1
XU$$4452 _582_/Q U$$4388/X _583_/Q U$$4468/B2 VGND VGND VPWR VPWR U$$4453/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_2 dadda_fa_2_49_2/A dadda_fa_2_49_2/B dadda_fa_2_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/A dadda_fa_3_49_3/A sky130_fd_sc_hd__fa_1
XFILLER_64_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4463 U$$4463/A U$$4463/B VGND VGND VPWR VPWR U$$4463/X sky130_fd_sc_hd__xor2_1
XFILLER_42_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4474 U$$4474/A1 U$$4388/X U$$4476/A1 U$$4480/B2 VGND VGND VPWR VPWR U$$4475/A
+ sky130_fd_sc_hd__a22o_1
XU$$4485 U$$4485/A U$$4485/B VGND VGND VPWR VPWR U$$4485/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_26_1 dadda_fa_5_26_1/A dadda_fa_5_26_1/B dadda_fa_5_26_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_27_0/B dadda_fa_7_26_0/A sky130_fd_sc_hd__fa_2
XU$$3740 U$$3740/A U$$3740/B VGND VGND VPWR VPWR U$$3740/X sky130_fd_sc_hd__xor2_1
XU$$3751 U$$3751/A1 U$$3785/A2 U$$3753/A1 U$$3785/B2 VGND VGND VPWR VPWR U$$3752/A
+ sky130_fd_sc_hd__a22o_1
XU$$4496 U$$934/A1 U$$4388/X U$$936/A1 U$$4496/B2 VGND VGND VPWR VPWR U$$4497/A sky130_fd_sc_hd__a22o_1
XU$$3762 U$$3762/A U$$3764/B VGND VGND VPWR VPWR U$$3762/X sky130_fd_sc_hd__xor2_1
XFILLER_25_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3773 U$$4456/B1 U$$3777/A2 U$$4323/A1 U$$3777/B2 VGND VGND VPWR VPWR U$$3774/A
+ sky130_fd_sc_hd__a22o_1
XU$$3784 U$$3784/A U$$3800/B VGND VGND VPWR VPWR U$$3784/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_19_0 dadda_fa_5_19_0/A dadda_fa_5_19_0/B dadda_fa_5_19_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_20_0/A dadda_fa_6_19_0/CIN sky130_fd_sc_hd__fa_2
XU$$3795 U$$3932/A1 U$$3795/A2 _597_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3796/A sky130_fd_sc_hd__a22o_1
XFILLER_64_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_100_1 dadda_fa_5_100_1/A dadda_fa_5_100_1/B dadda_fa_5_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_101_0/B dadda_fa_7_100_0/A sky130_fd_sc_hd__fa_2
XFILLER_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_4_122_0 dadda_ha_4_122_0/A U$$4108/X VGND VGND VPWR VPWR dadda_fa_5_123_1/CIN
+ dadda_ha_4_122_0/SUM sky130_fd_sc_hd__ha_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_556 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_38_2 U$$881/X U$$1014/X VGND VGND VPWR VPWR dadda_fa_2_39_5/A dadda_fa_3_38_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_102_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_96_0_1874 VGND VGND VPWR VPWR dadda_ha_1_96_0/A dadda_ha_1_96_0_1874/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_75_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_51_2 U$$907/X U$$1040/X U$$1173/X VGND VGND VPWR VPWR dadda_fa_2_52_1/A
+ dadda_fa_2_51_4/A sky130_fd_sc_hd__fa_1
XFILLER_84_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$906 U$$906/A1 U$$906/A2 U$$908/A1 U$$906/B2 VGND VGND VPWR VPWR U$$907/A sky130_fd_sc_hd__a22o_1
XFILLER_56_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$917 U$$917/A U$$958/A VGND VGND VPWR VPWR U$$917/X sky130_fd_sc_hd__xor2_1
XU$$928 U$$928/A1 U$$928/A2 U$$930/A1 U$$928/B2 VGND VGND VPWR VPWR U$$929/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_44_1 U$$494/X U$$627/X U$$760/X VGND VGND VPWR VPWR dadda_fa_2_45_2/CIN
+ dadda_fa_2_44_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_141_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$939 U$$939/A _629_/Q VGND VGND VPWR VPWR U$$939/X sky130_fd_sc_hd__xor2_1
XFILLER_43_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_21_0 input170/X dadda_fa_4_21_0/B dadda_fa_4_21_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_5_22_0/A dadda_fa_5_21_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_37_0 U$$81/X U$$214/X U$$347/X VGND VGND VPWR VPWR dadda_fa_2_38_4/CIN
+ dadda_fa_2_37_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_935 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_73_3 dadda_fa_3_73_3/A dadda_fa_3_73_3/B dadda_fa_3_73_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_1/B dadda_fa_4_73_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_692 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_66_2 dadda_fa_3_66_2/A dadda_fa_3_66_2/B dadda_fa_3_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_1/A dadda_fa_4_66_2/B sky130_fd_sc_hd__fa_1
XFILLER_120_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_59_1 dadda_fa_3_59_1/A dadda_fa_3_59_1/B dadda_fa_3_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_0/CIN dadda_fa_4_59_2/A sky130_fd_sc_hd__fa_1
XFILLER_78_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_36_0 dadda_fa_6_36_0/A dadda_fa_6_36_0/B dadda_fa_6_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_37_0/B dadda_fa_7_36_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3003 U$$3412/B1 U$$3005/A2 U$$3005/A1 U$$3005/B2 VGND VGND VPWR VPWR U$$3004/A
+ sky130_fd_sc_hd__a22o_1
XU$$3014 U$$3014/A VGND VGND VPWR VPWR U$$3014/Y sky130_fd_sc_hd__inv_1
XFILLER_74_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3025 U$$3025/A U$$3077/B VGND VGND VPWR VPWR U$$3025/X sky130_fd_sc_hd__xor2_1
XU$$3036 U$$3310/A1 U$$3046/A2 U$$3175/A1 U$$3046/B2 VGND VGND VPWR VPWR U$$3037/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2302 U$$2848/B1 U$$2302/A2 U$$658/B1 U$$2302/B2 VGND VGND VPWR VPWR U$$2303/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3047 U$$3047/A U$$3049/B VGND VGND VPWR VPWR U$$3047/X sky130_fd_sc_hd__xor2_1
XU$$3058 U$$42/B1 U$$3066/A2 U$$731/A1 U$$3066/B2 VGND VGND VPWR VPWR U$$3059/A sky130_fd_sc_hd__a22o_1
XU$$2313 U$$2313/A U$$2321/B VGND VGND VPWR VPWR U$$2313/X sky130_fd_sc_hd__xor2_1
XU$$2324 U$$954/A1 U$$2326/A2 U$$956/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2325/A sky130_fd_sc_hd__a22o_1
XU$$3069 U$$3069/A U$$3107/B VGND VGND VPWR VPWR U$$3069/X sky130_fd_sc_hd__xor2_1
XU$$2335 U$$2335/A1 U$$2367/A2 U$$2611/A1 U$$2367/B2 VGND VGND VPWR VPWR U$$2336/A
+ sky130_fd_sc_hd__a22o_1
XU$$1601 U$$2832/B1 U$$1607/A2 U$$2971/B1 U$$1607/B2 VGND VGND VPWR VPWR U$$1602/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2346 U$$2346/A U$$2366/B VGND VGND VPWR VPWR U$$2346/X sky130_fd_sc_hd__xor2_1
XU$$2357 U$$302/A1 U$$2387/A2 U$$2494/B1 U$$2387/B2 VGND VGND VPWR VPWR U$$2358/A
+ sky130_fd_sc_hd__a22o_1
XU$$1612 U$$1612/A U$$1636/B VGND VGND VPWR VPWR U$$1612/X sky130_fd_sc_hd__xor2_1
XU$$1623 U$$2991/B1 U$$1627/A2 U$$2858/A1 U$$1627/B2 VGND VGND VPWR VPWR U$$1624/A
+ sky130_fd_sc_hd__a22o_1
XU$$2368 U$$2368/A U$$2418/B VGND VGND VPWR VPWR U$$2368/X sky130_fd_sc_hd__xor2_1
XU$$2379 U$$4160/A1 U$$2435/A2 U$$4160/B1 U$$2435/B2 VGND VGND VPWR VPWR U$$2380/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1634 U$$1634/A U$$1636/B VGND VGND VPWR VPWR U$$1634/X sky130_fd_sc_hd__xor2_1
XU$$1645 _640_/Q VGND VGND VPWR VPWR U$$1647/B sky130_fd_sc_hd__inv_1
XFILLER_188_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1656 U$$971/A1 U$$1684/A2 U$$973/A1 U$$1684/B2 VGND VGND VPWR VPWR U$$1657/A sky130_fd_sc_hd__a22o_1
XU$$1667 U$$1667/A U$$1719/B VGND VGND VPWR VPWR U$$1667/X sky130_fd_sc_hd__xor2_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1678 U$$582/A1 U$$1718/A2 U$$582/B1 U$$1718/B2 VGND VGND VPWR VPWR U$$1679/A sky130_fd_sc_hd__a22o_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1689 U$$1689/A U$$1737/B VGND VGND VPWR VPWR U$$1689/X sky130_fd_sc_hd__xor2_1
XFILLER_202_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_309_ _439_/CLK _309_/D VGND VGND VPWR VPWR _309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_109_0 dadda_fa_7_109_0/A dadda_fa_7_109_0/B dadda_fa_7_109_0/CIN VGND
+ VGND VPWR VPWR _534_/D _405_/D sky130_fd_sc_hd__fa_1
XFILLER_162_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_61_1 dadda_fa_2_61_1/A dadda_fa_2_61_1/B dadda_fa_2_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_0/CIN dadda_fa_3_61_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater501 U$$3155/X VGND VGND VPWR VPWR U$$3283/A2 sky130_fd_sc_hd__buf_4
XFILLER_112_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$308 final_adder.U$$308/A final_adder.U$$308/B VGND VGND VPWR VPWR
+ final_adder.U$$346/B sky130_fd_sc_hd__and2_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater512 U$$2943/A2 VGND VGND VPWR VPWR U$$2915/A2 sky130_fd_sc_hd__buf_4
Xrepeater523 U$$392/A2 VGND VGND VPWR VPWR U$$350/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_54_0 dadda_fa_2_54_0/A dadda_fa_2_54_0/B dadda_fa_2_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_0/B dadda_fa_3_54_2/B sky130_fd_sc_hd__fa_2
Xrepeater534 U$$2744/X VGND VGND VPWR VPWR U$$2874/A2 sky130_fd_sc_hd__buf_6
XFILLER_84_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater545 U$$2524/A2 VGND VGND VPWR VPWR U$$2516/A2 sky130_fd_sc_hd__buf_4
Xrepeater556 U$$2451/A2 VGND VGND VPWR VPWR U$$2463/A2 sky130_fd_sc_hd__buf_6
Xrepeater567 U$$2135/A2 VGND VGND VPWR VPWR U$$2129/A2 sky130_fd_sc_hd__buf_4
XFILLER_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4260 U$$4260/A U$$4298/B VGND VGND VPWR VPWR U$$4260/X sky130_fd_sc_hd__xor2_1
Xrepeater578 U$$2038/A2 VGND VGND VPWR VPWR U$$2010/A2 sky130_fd_sc_hd__buf_6
XFILLER_81_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater589 U$$1907/A2 VGND VGND VPWR VPWR U$$1909/A2 sky130_fd_sc_hd__buf_6
XU$$4271 U$$4408/A1 U$$4297/A2 U$$4273/A1 U$$4297/B2 VGND VGND VPWR VPWR U$$4272/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4282 U$$4282/A U$$4322/B VGND VGND VPWR VPWR U$$4282/X sky130_fd_sc_hd__xor2_1
XU$$4293 U$$4293/A1 U$$4311/A2 _572_/Q U$$4311/B2 VGND VGND VPWR VPWR U$$4294/A sky130_fd_sc_hd__a22o_1
XU$$3570 U$$3844/A1 U$$3612/A2 _553_/Q U$$3612/B2 VGND VGND VPWR VPWR U$$3571/A sky130_fd_sc_hd__a22o_1
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3581 U$$3581/A U$$3609/B VGND VGND VPWR VPWR U$$3581/X sky130_fd_sc_hd__xor2_1
XU$$3592 U$$4003/A1 U$$3636/A2 U$$4140/B1 U$$3636/B2 VGND VGND VPWR VPWR U$$3593/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2880 U$$3014/A U$$2880/B VGND VGND VPWR VPWR U$$2880/X sky130_fd_sc_hd__and2_1
Xdadda_fa_5_8_0 U$$289/X U$$422/X U$$555/X VGND VGND VPWR VPWR dadda_fa_6_9_0/A dadda_fa_6_8_0/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_209_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2891 U$$3163/B1 U$$2943/A2 U$$3713/B1 U$$2943/B2 VGND VGND VPWR VPWR U$$2892/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4397_1777 VGND VGND VPWR VPWR U$$4397_1777/HI U$$4397/B sky130_fd_sc_hd__conb_1
XFILLER_88_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_83_2 dadda_fa_4_83_2/A dadda_fa_4_83_2/B dadda_fa_4_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/CIN dadda_fa_5_83_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_76_1 dadda_fa_4_76_1/A dadda_fa_4_76_1/B dadda_fa_4_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/B dadda_fa_5_76_1/B sky130_fd_sc_hd__fa_1
XFILLER_1_926 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_53_0 dadda_fa_7_53_0/A dadda_fa_7_53_0/B dadda_fa_7_53_0/CIN VGND VGND
+ VPWR VPWR _478_/D _349_/D sky130_fd_sc_hd__fa_1
XFILLER_103_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_69_0 dadda_fa_4_69_0/A dadda_fa_4_69_0/B dadda_fa_4_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/A dadda_fa_5_69_1/A sky130_fd_sc_hd__fa_1
XFILLER_130_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_660_ _660_/CLK _660_/D VGND VGND VPWR VPWR _660_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$703 U$$840/A1 U$$725/A2 U$$705/A1 U$$725/B2 VGND VGND VPWR VPWR U$$704/A sky130_fd_sc_hd__a22o_1
XFILLER_72_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$714 U$$714/A U$$766/B VGND VGND VPWR VPWR U$$714/X sky130_fd_sc_hd__xor2_1
XFILLER_1_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_591_ _596_/CLK _591_/D VGND VGND VPWR VPWR _591_/Q sky130_fd_sc_hd__dfxtp_1
XU$$725 U$$40/A1 U$$725/A2 U$$42/A1 U$$725/B2 VGND VGND VPWR VPWR U$$726/A sky130_fd_sc_hd__a22o_1
XFILLER_44_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$736 U$$736/A U$$748/B VGND VGND VPWR VPWR U$$736/X sky130_fd_sc_hd__xor2_1
XFILLER_17_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$747 U$$882/B1 U$$747/A2 U$$747/B1 U$$747/B2 VGND VGND VPWR VPWR U$$748/A sky130_fd_sc_hd__a22o_1
XFILLER_83_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$758 U$$758/A U$$804/B VGND VGND VPWR VPWR U$$758/X sky130_fd_sc_hd__xor2_1
XU$$769 U$$906/A1 U$$783/A2 U$$84/B1 U$$783/B2 VGND VGND VPWR VPWR U$$770/A sky130_fd_sc_hd__a22o_1
XFILLER_44_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1603 U$$3181/B1 VGND VGND VPWR VPWR U$$715/B1 sky130_fd_sc_hd__buf_6
XFILLER_153_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1614 U$$2494/B1 VGND VGND VPWR VPWR U$$989/A1 sky130_fd_sc_hd__buf_4
XANTENNA_8 _472_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1625 U$$4273/B1 VGND VGND VPWR VPWR U$$4136/B1 sky130_fd_sc_hd__buf_6
Xrepeater1636 _561_/Q VGND VGND VPWR VPWR U$$4273/A1 sky130_fd_sc_hd__buf_6
XFILLER_126_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1647 U$$22/A1 VGND VGND VPWR VPWR U$$20/B1 sky130_fd_sc_hd__buf_6
Xrepeater1658 U$$3717/B1 VGND VGND VPWR VPWR U$$840/B1 sky130_fd_sc_hd__buf_4
XFILLER_193_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1669 _557_/Q VGND VGND VPWR VPWR U$$2893/B1 sky130_fd_sc_hd__buf_4
XFILLER_3_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_71_0 dadda_fa_3_71_0/A dadda_fa_3_71_0/B dadda_fa_3_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_0/B dadda_fa_4_71_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2110 U$$2110/A U$$2110/B VGND VGND VPWR VPWR U$$2110/X sky130_fd_sc_hd__xor2_1
XFILLER_63_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_100_0 dadda_fa_4_100_0/A dadda_fa_4_100_0/B dadda_fa_4_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/A dadda_fa_5_100_1/A sky130_fd_sc_hd__fa_1
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2121 U$$3626/B1 U$$2135/A2 U$$3493/A1 U$$2135/B2 VGND VGND VPWR VPWR U$$2122/A
+ sky130_fd_sc_hd__a22o_1
XU$$2132 U$$2132/A U$$2136/B VGND VGND VPWR VPWR U$$2132/X sky130_fd_sc_hd__xor2_1
XFILLER_63_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2143 U$$2963/B1 U$$2145/A2 U$$2830/A1 U$$2145/B2 VGND VGND VPWR VPWR U$$2144/A
+ sky130_fd_sc_hd__a22o_1
XU$$2154 U$$2154/A U$$2191/A VGND VGND VPWR VPWR U$$2154/X sky130_fd_sc_hd__xor2_1
XFILLER_23_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1420 U$$596/B1 U$$1458/A2 U$$463/A1 U$$1458/B2 VGND VGND VPWR VPWR U$$1421/A sky130_fd_sc_hd__a22o_1
XU$$2165 U$$2848/B1 U$$2169/A2 U$$2715/A1 U$$2169/B2 VGND VGND VPWR VPWR U$$2166/A
+ sky130_fd_sc_hd__a22o_1
XU$$2176 U$$2176/A U$$2186/B VGND VGND VPWR VPWR U$$2176/X sky130_fd_sc_hd__xor2_1
XU$$1431 U$$1431/A U$$1479/B VGND VGND VPWR VPWR U$$1431/X sky130_fd_sc_hd__xor2_1
XU$$1442 U$$3221/B1 U$$1442/A2 U$$74/A1 U$$1442/B2 VGND VGND VPWR VPWR U$$1443/A sky130_fd_sc_hd__a22o_1
XU$$2187 U$$2459/B1 U$$2189/A2 U$$956/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2188/A
+ sky130_fd_sc_hd__a22o_1
XU$$1453 U$$1453/A U$$1479/B VGND VGND VPWR VPWR U$$1453/X sky130_fd_sc_hd__xor2_1
XU$$2198 U$$2198/A1 U$$2248/A2 U$$2611/A1 U$$2248/B2 VGND VGND VPWR VPWR U$$2199/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1464 U$$94/A1 U$$1474/A2 U$$2971/B1 U$$1474/B2 VGND VGND VPWR VPWR U$$1465/A sky130_fd_sc_hd__a22o_1
XFILLER_96_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1475 U$$1475/A U$$1475/B VGND VGND VPWR VPWR U$$1475/X sky130_fd_sc_hd__xor2_1
XFILLER_194_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1486 U$$251/B1 U$$1486/A2 U$$2858/A1 U$$1486/B2 VGND VGND VPWR VPWR U$$1487/A
+ sky130_fd_sc_hd__a22o_1
XU$$1497 U$$1497/A U$$1501/B VGND VGND VPWR VPWR U$$1497/X sky130_fd_sc_hd__xor2_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_93_1 dadda_fa_5_93_1/A dadda_fa_5_93_1/B dadda_fa_5_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_94_0/B dadda_fa_7_93_0/A sky130_fd_sc_hd__fa_1
XFILLER_117_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_580 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_86_0 dadda_fa_5_86_0/A dadda_fa_5_86_0/B dadda_fa_5_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_87_0/A dadda_fa_6_86_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_190_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_78_7 U$$4020/X U$$4153/X U$$4286/X VGND VGND VPWR VPWR dadda_fa_2_79_2/CIN
+ dadda_fa_2_78_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$105 _529_/Q _401_/Q VGND VGND VPWR VPWR final_adder.U$$233/B1 final_adder.U$$727/A
+ sky130_fd_sc_hd__ha_2
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_1028 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$116 _540_/Q _412_/Q VGND VGND VPWR VPWR final_adder.U$$611/B1 final_adder.U$$738/A
+ sky130_fd_sc_hd__ha_2
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$127 _551_/Q _423_/Q VGND VGND VPWR VPWR final_adder.U$$127/COUT final_adder.U$$749/A
+ sky130_fd_sc_hd__ha_1
XFILLER_57_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$138 final_adder.U$$633/A final_adder.U$$632/A VGND VGND VPWR VPWR
+ final_adder.U$$260/A sky130_fd_sc_hd__and2_1
XFILLER_211_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$149 final_adder.U$$643/A final_adder.U$$515/B1 final_adder.U$$149/B1
+ VGND VGND VPWR VPWR final_adder.U$$149/X sky130_fd_sc_hd__a21o_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater386 U$$999/A2 VGND VGND VPWR VPWR U$$979/A2 sky130_fd_sc_hd__buf_4
XFILLER_38_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater397 U$$924/A2 VGND VGND VPWR VPWR U$$896/A2 sky130_fd_sc_hd__buf_4
XU$$4090 U$$4090/A U$$4096/B VGND VGND VPWR VPWR U$$4090/X sky130_fd_sc_hd__xor2_1
XFILLER_38_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_868 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_102_2 dadda_fa_3_102_2/A dadda_fa_3_102_2/B dadda_fa_3_102_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_103_1/A dadda_fa_4_102_2/B sky130_fd_sc_hd__fa_1
XFILLER_134_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 b[42] VGND VGND VPWR VPWR _594_/D sky130_fd_sc_hd__clkbuf_1
Xinput112 b[52] VGND VGND VPWR VPWR _604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput123 b[62] VGND VGND VPWR VPWR _614_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput134 c[104] VGND VGND VPWR VPWR input134/X sky130_fd_sc_hd__buf_2
XTAP_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput145 c[114] VGND VGND VPWR VPWR input145/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_66_5 U$$2134/X U$$2267/X U$$2400/X VGND VGND VPWR VPWR dadda_fa_1_67_7/A
+ dadda_fa_2_66_0/A sky130_fd_sc_hd__fa_2
Xinput156 c[124] VGND VGND VPWR VPWR input156/X sky130_fd_sc_hd__clkbuf_1
XTAP_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_116_0 dadda_fa_6_116_0/A dadda_fa_6_116_0/B dadda_fa_6_116_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_117_0/B dadda_fa_7_116_0/CIN sky130_fd_sc_hd__fa_1
Xinput167 c[19] VGND VGND VPWR VPWR input167/X sky130_fd_sc_hd__buf_2
XTAP_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput178 c[29] VGND VGND VPWR VPWR input178/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1041 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 c[39] VGND VGND VPWR VPWR input189/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$650 final_adder.U$$650/A final_adder.U$$650/B VGND VGND VPWR VPWR
+ _196_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$661 final_adder.U$$661/A final_adder.U$$661/B VGND VGND VPWR VPWR
+ _207_/D sky130_fd_sc_hd__xor2_1
XTAP_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$500 U$$500/A U$$500/B VGND VGND VPWR VPWR U$$500/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$672 final_adder.U$$672/A final_adder.U$$672/B VGND VGND VPWR VPWR
+ _218_/D sky130_fd_sc_hd__xor2_1
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$511 U$$648/A1 U$$517/A2 U$$648/B1 U$$517/B2 VGND VGND VPWR VPWR U$$512/A sky130_fd_sc_hd__a22o_1
X_643_ _648_/CLK _643_/D VGND VGND VPWR VPWR _643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_36_3 dadda_fa_3_36_3/A dadda_fa_3_36_3/B dadda_fa_3_36_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_1/B dadda_fa_4_36_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$683 final_adder.U$$683/A final_adder.U$$683/B VGND VGND VPWR VPWR
+ _229_/D sky130_fd_sc_hd__xor2_1
XTAP_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$522 U$$522/A U$$547/A VGND VGND VPWR VPWR U$$522/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$694 final_adder.U$$694/A final_adder.U$$694/B VGND VGND VPWR VPWR
+ _240_/D sky130_fd_sc_hd__xor2_1
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$533 U$$805/B1 U$$415/X U$$944/B1 U$$416/X VGND VGND VPWR VPWR U$$534/A sky130_fd_sc_hd__a22o_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$544 U$$544/A U$$547/A VGND VGND VPWR VPWR U$$544/X sky130_fd_sc_hd__xor2_1
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$555 U$$555/A U$$627/B VGND VGND VPWR VPWR U$$555/X sky130_fd_sc_hd__xor2_1
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_574_ _575_/CLK _574_/D VGND VGND VPWR VPWR _574_/Q sky130_fd_sc_hd__dfxtp_4
XU$$566 U$$840/A1 U$$574/A2 U$$705/A1 U$$574/B2 VGND VGND VPWR VPWR U$$567/A sky130_fd_sc_hd__a22o_1
XFILLER_17_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_29_2 dadda_fa_3_29_2/A dadda_fa_3_29_2/B dadda_fa_3_29_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_30_1/A dadda_fa_4_29_2/B sky130_fd_sc_hd__fa_1
XU$$577 U$$577/A U$$613/B VGND VGND VPWR VPWR U$$577/X sky130_fd_sc_hd__xor2_1
XU$$588 U$$40/A1 U$$622/A2 U$$42/A1 U$$622/B2 VGND VGND VPWR VPWR U$$589/A sky130_fd_sc_hd__a22o_1
XU$$599 U$$599/A U$$627/B VGND VGND VPWR VPWR U$$599/X sky130_fd_sc_hd__xor2_1
XFILLER_72_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1400 U$$3646/A1 VGND VGND VPWR VPWR U$$3372/A1 sky130_fd_sc_hd__buf_6
Xrepeater1411 U$$900/B1 VGND VGND VPWR VPWR U$$80/A1 sky130_fd_sc_hd__buf_4
Xrepeater1422 U$$4051/A1 VGND VGND VPWR VPWR U$$3229/A1 sky130_fd_sc_hd__buf_4
Xrepeater1433 U$$4323/A1 VGND VGND VPWR VPWR U$$4186/A1 sky130_fd_sc_hd__buf_6
XFILLER_67_1025 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1444 U$$2947/B1 VGND VGND VPWR VPWR U$$894/A1 sky130_fd_sc_hd__buf_6
Xrepeater1455 _583_/Q VGND VGND VPWR VPWR U$$3221/A1 sky130_fd_sc_hd__buf_4
XFILLER_141_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1466 _582_/Q VGND VGND VPWR VPWR U$$4176/B1 sky130_fd_sc_hd__buf_4
XFILLER_141_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1477 U$$201/A1 VGND VGND VPWR VPWR U$$64/A1 sky130_fd_sc_hd__buf_4
XFILLER_99_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1488 U$$3624/A1 VGND VGND VPWR VPWR U$$3896/B1 sky130_fd_sc_hd__buf_8
Xrepeater1499 _578_/Q VGND VGND VPWR VPWR U$$4444/A1 sky130_fd_sc_hd__buf_8
XFILLER_80_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_31_2 U$$867/X U$$1000/X U$$1133/X VGND VGND VPWR VPWR dadda_fa_3_32_1/B
+ dadda_fa_3_31_3/B sky130_fd_sc_hd__fa_1
XFILLER_39_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1250 U$$1250/A U$$1296/B VGND VGND VPWR VPWR U$$1250/X sky130_fd_sc_hd__xor2_1
XFILLER_189_971 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1261 U$$302/A1 U$$1323/A2 U$$989/A1 U$$1323/B2 VGND VGND VPWR VPWR U$$1262/A sky130_fd_sc_hd__a22o_1
XFILLER_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1272 U$$1272/A U$$1280/B VGND VGND VPWR VPWR U$$1272/X sky130_fd_sc_hd__xor2_1
XFILLER_176_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1283 U$$733/B1 U$$1291/A2 U$$600/A1 U$$1291/B2 VGND VGND VPWR VPWR U$$1284/A sky130_fd_sc_hd__a22o_1
XFILLER_176_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1294 U$$1294/A U$$1332/B VGND VGND VPWR VPWR U$$1294/X sky130_fd_sc_hd__xor2_1
XFILLER_191_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_83_5 U$$3365/X U$$3498/X U$$3631/X VGND VGND VPWR VPWR dadda_fa_2_84_3/B
+ dadda_fa_2_83_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_76_4 U$$3085/X U$$3218/X U$$3351/X VGND VGND VPWR VPWR dadda_fa_2_77_1/CIN
+ dadda_fa_2_76_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_3 U$$3603/X U$$3736/X U$$3869/X VGND VGND VPWR VPWR dadda_fa_2_70_1/B
+ dadda_fa_2_69_4/B sky130_fd_sc_hd__fa_1
XFILLER_97_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_46_2 dadda_fa_4_46_2/A dadda_fa_4_46_2/B dadda_fa_4_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/CIN dadda_fa_5_46_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_39_1 dadda_fa_4_39_1/A dadda_fa_4_39_1/B dadda_fa_4_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/B dadda_fa_5_39_1/B sky130_fd_sc_hd__fa_1
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_7_16_0 dadda_fa_7_16_0/A dadda_fa_7_16_0/B dadda_fa_7_16_0/CIN VGND VGND
+ VPWR VPWR _441_/D _312_/D sky130_fd_sc_hd__fa_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_228 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_239 _192_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_290_ _615_/CLK _290_/D VGND VGND VPWR VPWR _290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_58_3 U$$1320/X U$$1453/X VGND VGND VPWR VPWR dadda_fa_1_59_7/CIN dadda_fa_2_58_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_71_3 U$$1745/X U$$1878/X U$$2011/X VGND VGND VPWR VPWR dadda_fa_1_72_7/CIN
+ dadda_fa_2_71_0/A sky130_fd_sc_hd__fa_1
XTAP_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_64_2 U$$933/X U$$1066/X U$$1199/X VGND VGND VPWR VPWR dadda_fa_1_65_6/A
+ dadda_fa_1_64_8/A sky130_fd_sc_hd__fa_1
XFILLER_7_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_41_1 dadda_fa_3_41_1/A dadda_fa_3_41_1/B dadda_fa_3_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_0/CIN dadda_fa_4_41_2/A sky130_fd_sc_hd__fa_1
XTAP_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_57_1 U$$520/X U$$653/X U$$786/X VGND VGND VPWR VPWR dadda_fa_1_58_7/B
+ dadda_fa_1_57_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_188_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_34_0 dadda_fa_3_34_0/A dadda_fa_3_34_0/B dadda_fa_3_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_0/B dadda_fa_4_34_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$491 final_adder.U$$314/B final_adder.U$$738/B final_adder.U$$245/X
+ VGND VGND VPWR VPWR final_adder.U$$740/B sky130_fd_sc_hd__a21o_1
XU$$330 U$$330/A1 U$$398/A2 U$$58/A1 U$$398/B2 VGND VGND VPWR VPWR U$$331/A sky130_fd_sc_hd__a22o_1
X_626_ _626_/CLK _626_/D VGND VGND VPWR VPWR _626_/Q sky130_fd_sc_hd__dfxtp_2
XU$$341 U$$341/A U$$351/B VGND VGND VPWR VPWR U$$341/X sky130_fd_sc_hd__xor2_1
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$352 U$$624/B1 U$$398/A2 U$$491/A1 U$$398/B2 VGND VGND VPWR VPWR U$$353/A sky130_fd_sc_hd__a22o_1
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$363 U$$363/A U$$410/A VGND VGND VPWR VPWR U$$363/X sky130_fd_sc_hd__xor2_1
XFILLER_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$374 U$$648/A1 U$$384/A2 U$$648/B1 U$$384/B2 VGND VGND VPWR VPWR U$$375/A sky130_fd_sc_hd__a22o_1
XFILLER_45_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$385 U$$385/A U$$393/B VGND VGND VPWR VPWR U$$385/X sky130_fd_sc_hd__xor2_1
XFILLER_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_557_ _559_/CLK _557_/D VGND VGND VPWR VPWR _557_/Q sky130_fd_sc_hd__dfxtp_4
XU$$396 U$$805/B1 U$$398/A2 U$$944/B1 U$$398/B2 VGND VGND VPWR VPWR U$$397/A sky130_fd_sc_hd__a22o_1
XFILLER_33_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_488_ _488_/CLK _488_/D VGND VGND VPWR VPWR _488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_93_4 U$$4449/X input249/X dadda_fa_2_93_4/CIN VGND VGND VPWR VPWR dadda_fa_3_94_1/CIN
+ dadda_fa_3_93_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1230 U$$2866/A1 VGND VGND VPWR VPWR U$$3412/B1 sky130_fd_sc_hd__buf_6
XFILLER_59_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1241 U$$2586/B1 VGND VGND VPWR VPWR U$$944/A1 sky130_fd_sc_hd__buf_6
Xrepeater1252 U$$940/B1 VGND VGND VPWR VPWR U$$4504/A1 sky130_fd_sc_hd__buf_8
Xrepeater1263 U$$3132/A1 VGND VGND VPWR VPWR U$$2858/A1 sky130_fd_sc_hd__buf_6
XFILLER_5_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_86_3 dadda_fa_2_86_3/A dadda_fa_2_86_3/B dadda_fa_2_86_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_1/B dadda_fa_3_86_3/B sky130_fd_sc_hd__fa_1
Xrepeater1274 _605_/Q VGND VGND VPWR VPWR U$$2991/A1 sky130_fd_sc_hd__buf_4
Xrepeater1285 U$$4494/B1 VGND VGND VPWR VPWR U$$934/A1 sky130_fd_sc_hd__buf_4
XFILLER_114_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1296 U$$3807/B1 VGND VGND VPWR VPWR U$$4355/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_79_2 dadda_fa_2_79_2/A dadda_fa_2_79_2/B dadda_fa_2_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/A dadda_fa_3_79_3/A sky130_fd_sc_hd__fa_1
XFILLER_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_56_1 dadda_fa_5_56_1/A dadda_fa_5_56_1/B dadda_fa_5_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_57_0/B dadda_fa_7_56_0/A sky130_fd_sc_hd__fa_1
XFILLER_113_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_952 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_49_0 dadda_fa_5_49_0/A dadda_fa_5_49_0/B dadda_fa_5_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_50_0/A dadda_fa_6_49_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_2_23_0 U$$53/X U$$186/X VGND VGND VPWR VPWR dadda_fa_3_24_3/B dadda_fa_4_23_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_95_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_102_1 U$$3004/X U$$3137/X U$$3270/X VGND VGND VPWR VPWR dadda_fa_3_103_2/B
+ dadda_fa_3_102_3/B sky130_fd_sc_hd__fa_1
XFILLER_63_582 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1080 U$$1080/A U$$1095/A VGND VGND VPWR VPWR U$$1080/X sky130_fd_sc_hd__xor2_1
XFILLER_17_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1091 U$$954/A1 U$$1093/A2 U$$956/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1092/A sky130_fd_sc_hd__a22o_1
XFILLER_32_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_123_0 U$$4109/Y U$$4243/X U$$4376/X VGND VGND VPWR VPWR dadda_fa_6_124_0/A
+ dadda_fa_6_123_0/CIN sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_30_clk _479_/CLK VGND VGND VPWR VPWR _476_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_81_2 U$$2031/X U$$2164/X U$$2297/X VGND VGND VPWR VPWR dadda_fa_2_82_1/CIN
+ dadda_fa_2_81_4/B sky130_fd_sc_hd__fa_1
XFILLER_137_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_74_1 U$$2150/X U$$2283/X U$$2416/X VGND VGND VPWR VPWR dadda_fa_2_75_0/CIN
+ dadda_fa_2_74_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_51_0 dadda_fa_4_51_0/A dadda_fa_4_51_0/B dadda_fa_4_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/A dadda_fa_5_51_1/A sky130_fd_sc_hd__fa_1
XFILLER_58_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_97_clk _634_/CLK VGND VGND VPWR VPWR _494_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_1_67_0 U$$2535/X U$$2668/X U$$2801/X VGND VGND VPWR VPWR dadda_fa_2_68_0/B
+ dadda_fa_2_67_3/B sky130_fd_sc_hd__fa_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2709 U$$3942/A1 U$$2607/X U$$4218/A1 U$$2608/X VGND VGND VPWR VPWR U$$2710/A sky130_fd_sc_hd__a22o_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_411_ _648_/CLK _411_/D VGND VGND VPWR VPWR _411_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_342_ _343_/CLK _342_/D VGND VGND VPWR VPWR _342_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_273_ _521_/CLK _273_/D VGND VGND VPWR VPWR _273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk _432_/CLK VGND VGND VPWR VPWR _431_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_808 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_96_2 dadda_fa_3_96_2/A dadda_fa_3_96_2/B dadda_fa_3_96_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_1/A dadda_fa_4_96_2/B sky130_fd_sc_hd__fa_1
XFILLER_68_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_89_1 dadda_fa_3_89_1/A dadda_fa_3_89_1/B dadda_fa_3_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_0/CIN dadda_fa_4_89_2/A sky130_fd_sc_hd__fa_1
XFILLER_120_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_66_0 dadda_fa_6_66_0/A dadda_fa_6_66_0/B dadda_fa_6_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_67_0/B dadda_fa_7_66_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_190_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_88_clk _628_/CLK VGND VGND VPWR VPWR _542_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater908 U$$4350/B VGND VGND VPWR VPWR U$$4348/B sky130_fd_sc_hd__buf_6
Xrepeater919 U$$4203/B VGND VGND VPWR VPWR U$$4247/A sky130_fd_sc_hd__buf_4
XFILLER_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3900 U$$4035/B1 U$$3958/A2 U$$4176/A1 U$$3958/B2 VGND VGND VPWR VPWR U$$3901/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3911 U$$3911/A U$$3933/B VGND VGND VPWR VPWR U$$3911/X sky130_fd_sc_hd__xor2_1
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_118_1 U$$4100/X U$$4233/X U$$4366/X VGND VGND VPWR VPWR dadda_fa_5_119_0/CIN
+ dadda_fa_5_118_1/B sky130_fd_sc_hd__fa_1
XFILLER_76_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3922 U$$4194/B1 U$$3932/A2 _592_/Q U$$3932/B2 VGND VGND VPWR VPWR U$$3923/A sky130_fd_sc_hd__a22o_1
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3933 U$$3933/A U$$3933/B VGND VGND VPWR VPWR U$$3933/X sky130_fd_sc_hd__xor2_1
XFILLER_40_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3944 U$$4218/A1 U$$3968/A2 U$$4355/B1 U$$3968/B2 VGND VGND VPWR VPWR U$$3945/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3955 U$$3955/A U$$3973/A VGND VGND VPWR VPWR U$$3955/X sky130_fd_sc_hd__xor2_1
XU$$3966 U$$4238/B1 U$$3970/A2 U$$4105/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3967/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3977 U$$3975/Y _674_/Q _673_/Q U$$3976/X U$$3973/Y VGND VGND VPWR VPWR U$$3977/X
+ sky130_fd_sc_hd__a32o_2
XU$$3988 U$$3988/A U$$3994/B VGND VGND VPWR VPWR U$$3988/X sky130_fd_sc_hd__xor2_1
XU$$160 U$$160/A U$$190/B VGND VGND VPWR VPWR U$$160/X sky130_fd_sc_hd__xor2_1
X_609_ _615_/CLK _609_/D VGND VGND VPWR VPWR _609_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3999 U$$4273/A1 U$$4035/A2 U$$4136/B1 U$$4081/B2 VGND VGND VPWR VPWR U$$4000/A
+ sky130_fd_sc_hd__a22o_1
XU$$171 U$$34/A1 U$$195/A2 U$$36/A1 U$$195/B2 VGND VGND VPWR VPWR U$$172/A sky130_fd_sc_hd__a22o_1
XU$$182 U$$182/A U$$216/B VGND VGND VPWR VPWR U$$182/X sky130_fd_sc_hd__xor2_1
XFILLER_33_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$193 U$$330/A1 U$$195/A2 U$$58/A1 U$$195/B2 VGND VGND VPWR VPWR U$$194/A sky130_fd_sc_hd__a22o_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_755 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_12_clk _616_/CLK VGND VGND VPWR VPWR _455_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_203_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_91_1 U$$3514/X U$$3647/X U$$3780/X VGND VGND VPWR VPWR dadda_fa_3_92_0/CIN
+ dadda_fa_3_91_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1060 U$$2039/B VGND VGND VPWR VPWR U$$2011/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_84_0 U$$4032/X U$$4165/X U$$4298/X VGND VGND VPWR VPWR dadda_fa_3_85_0/B
+ dadda_fa_3_84_2/B sky130_fd_sc_hd__fa_1
XFILLER_173_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput257 _168_/Q VGND VGND VPWR VPWR o[0] sky130_fd_sc_hd__buf_2
Xrepeater1071 U$$1916/B VGND VGND VPWR VPWR U$$1917/A sky130_fd_sc_hd__buf_6
Xoutput268 _178_/Q VGND VGND VPWR VPWR o[10] sky130_fd_sc_hd__buf_2
XFILLER_142_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1082 _641_/Q VGND VGND VPWR VPWR U$$1780/A sky130_fd_sc_hd__buf_6
Xoutput279 _179_/Q VGND VGND VPWR VPWR o[11] sky130_fd_sc_hd__buf_2
Xrepeater1093 U$$1475/B VGND VGND VPWR VPWR U$$1459/B sky130_fd_sc_hd__buf_6
XFILLER_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_60_7 dadda_fa_1_60_7/A dadda_fa_1_60_7/B dadda_fa_1_60_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_61_2/CIN dadda_fa_2_60_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_6 U$$2773/X U$$2906/X U$$3039/X VGND VGND VPWR VPWR dadda_fa_2_54_2/B
+ dadda_fa_2_53_5/B sky130_fd_sc_hd__fa_1
XFILLER_28_549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_46_5 U$$2094/X U$$2227/X U$$2360/X VGND VGND VPWR VPWR dadda_fa_2_47_3/B
+ dadda_fa_2_46_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_167_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_5_0 dadda_fa_7_5_0/A dadda_fa_7_5_0/B dadda_fa_7_5_0/CIN VGND VGND VPWR
+ VPWR _430_/D _301_/D sky130_fd_sc_hd__fa_1
XFILLER_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1011 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_83_0 dadda_fa_7_83_0/A dadda_fa_7_83_0/B dadda_fa_7_83_0/CIN VGND VGND
+ VPWR VPWR _508_/D _379_/D sky130_fd_sc_hd__fa_1
XFILLER_137_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_99_0 dadda_fa_4_99_0/A dadda_fa_4_99_0/B dadda_fa_4_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/A dadda_fa_5_99_1/A sky130_fd_sc_hd__fa_1
XFILLER_30_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1099 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3207 U$$4027/B1 U$$3285/A2 U$$467/B1 U$$3285/B2 VGND VGND VPWR VPWR U$$3208/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3218 U$$3218/A U$$3218/B VGND VGND VPWR VPWR U$$3218/X sky130_fd_sc_hd__xor2_1
XFILLER_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3229 U$$3229/A1 U$$3231/A2 U$$628/A1 U$$3231/B2 VGND VGND VPWR VPWR U$$3230/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2506 U$$2641/B1 U$$2550/A2 U$$2508/A1 U$$2550/B2 VGND VGND VPWR VPWR U$$2507/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2517 U$$2517/A U$$2517/B VGND VGND VPWR VPWR U$$2517/X sky130_fd_sc_hd__xor2_1
XU$$2528 U$$4035/A1 U$$2530/A2 U$$4035/B1 U$$2530/B2 VGND VGND VPWR VPWR U$$2529/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2539 U$$2539/A U$$2567/B VGND VGND VPWR VPWR U$$2539/X sky130_fd_sc_hd__xor2_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1805 U$$2077/B1 U$$1843/A2 U$$4410/A1 U$$1843/B2 VGND VGND VPWR VPWR U$$1806/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1816 U$$1816/A U$$1874/B VGND VGND VPWR VPWR U$$1816/X sky130_fd_sc_hd__xor2_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1827 U$$866/B1 U$$1855/A2 U$$2786/B1 U$$1855/B2 VGND VGND VPWR VPWR U$$1828/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1838 U$$1838/A U$$1844/B VGND VGND VPWR VPWR U$$1838/X sky130_fd_sc_hd__xor2_1
XFILLER_15_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1849 U$$68/A1 U$$1851/A2 U$$3358/A1 U$$1851/B2 VGND VGND VPWR VPWR U$$1850/A sky130_fd_sc_hd__a22o_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ _454_/CLK _325_/D VGND VGND VPWR VPWR _325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_256_ _519_/CLK _256_/D VGND VGND VPWR VPWR _256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_187_ _189_/CLK _187_/D VGND VGND VPWR VPWR _187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_896 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_63_5 dadda_fa_2_63_5/A dadda_fa_2_63_5/B dadda_fa_2_63_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_2/A dadda_fa_4_63_0/A sky130_fd_sc_hd__fa_2
XFILLER_85_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater705 U$$3910/B2 VGND VGND VPWR VPWR U$$3874/B2 sky130_fd_sc_hd__buf_4
Xrepeater716 U$$3805/B2 VGND VGND VPWR VPWR U$$3823/B2 sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_1_clk _442_/CLK VGND VGND VPWR VPWR _441_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater727 U$$3430/X VGND VGND VPWR VPWR U$$3497/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_56_4 dadda_fa_2_56_4/A dadda_fa_2_56_4/B dadda_fa_2_56_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/CIN dadda_fa_3_56_3/CIN sky130_fd_sc_hd__fa_1
XU$$4420 _566_/Q U$$4388/X _567_/Q U$$4454/B2 VGND VGND VPWR VPWR U$$4421/A sky130_fd_sc_hd__a22o_1
XFILLER_38_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater738 U$$3408/B2 VGND VGND VPWR VPWR U$$3378/B2 sky130_fd_sc_hd__buf_6
XFILLER_133_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater749 U$$3156/X VGND VGND VPWR VPWR U$$3283/B2 sky130_fd_sc_hd__buf_4
XU$$4431 U$$4431/A U$$4431/B VGND VGND VPWR VPWR U$$4431/X sky130_fd_sc_hd__xor2_1
XU$$4442 U$$4442/A1 U$$4388/X U$$4444/A1 U$$4454/B2 VGND VGND VPWR VPWR U$$4443/A
+ sky130_fd_sc_hd__a22o_1
XU$$4453 U$$4453/A U$$4453/B VGND VGND VPWR VPWR U$$4453/X sky130_fd_sc_hd__xor2_1
XFILLER_93_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4464 U$$4464/A1 U$$4388/X U$$4466/A1 U$$4468/B2 VGND VGND VPWR VPWR U$$4465/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_3 dadda_fa_2_49_3/A dadda_fa_2_49_3/B dadda_fa_2_49_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/B dadda_fa_3_49_3/B sky130_fd_sc_hd__fa_1
XFILLER_42_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3730 U$$3730/A U$$3832/B VGND VGND VPWR VPWR U$$3730/X sky130_fd_sc_hd__xor2_1
XFILLER_64_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4475 U$$4475/A U$$4475/B VGND VGND VPWR VPWR U$$4475/X sky130_fd_sc_hd__xor2_1
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4486 U$$4486/A1 U$$4388/X U$$926/A1 U$$4496/B2 VGND VGND VPWR VPWR U$$4487/A sky130_fd_sc_hd__a22o_1
XU$$3741 U$$3876/B1 U$$3743/A2 U$$3741/B1 U$$3743/B2 VGND VGND VPWR VPWR U$$3742/A
+ sky130_fd_sc_hd__a22o_1
XU$$3752 U$$3752/A U$$3760/B VGND VGND VPWR VPWR U$$3752/X sky130_fd_sc_hd__xor2_1
XU$$4497 U$$4497/A U$$4497/B VGND VGND VPWR VPWR U$$4497/X sky130_fd_sc_hd__xor2_1
XFILLER_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3763 U$$4448/A1 U$$3777/A2 U$$4176/A1 U$$3777/B2 VGND VGND VPWR VPWR U$$3764/A
+ sky130_fd_sc_hd__a22o_1
XU$$3774 U$$3774/A _671_/Q VGND VGND VPWR VPWR U$$3774/X sky130_fd_sc_hd__xor2_1
XU$$3785 U$$4194/B1 U$$3785/A2 U$$4061/A1 U$$3785/B2 VGND VGND VPWR VPWR U$$3786/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_19_1 dadda_fa_5_19_1/A dadda_fa_5_19_1/B dadda_fa_5_19_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_20_0/B dadda_fa_7_19_0/A sky130_fd_sc_hd__fa_2
XU$$3796 U$$3796/A U$$3800/B VGND VGND VPWR VPWR U$$3796/X sky130_fd_sc_hd__xor2_1
XFILLER_127_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_922 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_51_3 U$$1306/X U$$1439/X U$$1572/X VGND VGND VPWR VPWR dadda_fa_2_52_1/B
+ dadda_fa_2_51_4/B sky130_fd_sc_hd__fa_1
XU$$907 U$$907/A U$$907/B VGND VGND VPWR VPWR U$$907/X sky130_fd_sc_hd__xor2_1
XU$$918 U$$96/A1 U$$948/A2 U$$918/B1 U$$948/B2 VGND VGND VPWR VPWR U$$919/A sky130_fd_sc_hd__a22o_1
XU$$929 U$$929/A U$$929/B VGND VGND VPWR VPWR U$$929/X sky130_fd_sc_hd__xor2_1
XFILLER_56_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_44_2 U$$893/X U$$1026/X U$$1159/X VGND VGND VPWR VPWR dadda_fa_2_45_3/A
+ dadda_fa_2_44_5/A sky130_fd_sc_hd__fa_1
XFILLER_141_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_21_1 dadda_fa_4_21_1/A dadda_fa_4_21_1/B dadda_fa_4_21_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_22_0/B dadda_fa_5_21_1/B sky130_fd_sc_hd__fa_1
XFILLER_169_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_14_0 U$$301/X U$$434/X U$$567/X VGND VGND VPWR VPWR dadda_fa_5_15_0/A
+ dadda_fa_5_14_1/A sky130_fd_sc_hd__fa_1
XFILLER_197_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_66_3 dadda_fa_3_66_3/A dadda_fa_3_66_3/B dadda_fa_3_66_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_1/B dadda_fa_4_66_2/CIN sky130_fd_sc_hd__fa_1
XU$$4415_1786 VGND VGND VPWR VPWR U$$4415_1786/HI U$$4415/B sky130_fd_sc_hd__conb_1
Xdadda_fa_3_59_2 dadda_fa_3_59_2/A dadda_fa_3_59_2/B dadda_fa_3_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_1/A dadda_fa_4_59_2/B sky130_fd_sc_hd__fa_1
XFILLER_120_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3004 U$$3004/A U$$3008/B VGND VGND VPWR VPWR U$$3004/X sky130_fd_sc_hd__xor2_1
XU$$3015 _660_/Q VGND VGND VPWR VPWR U$$3017/B sky130_fd_sc_hd__inv_1
XFILLER_101_590 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_29_0 dadda_fa_6_29_0/A dadda_fa_6_29_0/B dadda_fa_6_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_30_0/B dadda_fa_7_29_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_806 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3026 U$$3437/A1 U$$3054/A2 U$$3163/B1 U$$3054/B2 VGND VGND VPWR VPWR U$$3027/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3037 U$$3037/A U$$3049/B VGND VGND VPWR VPWR U$$3037/X sky130_fd_sc_hd__xor2_1
XFILLER_74_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2303 U$$2303/A U$$2303/B VGND VGND VPWR VPWR U$$2303/X sky130_fd_sc_hd__xor2_1
XU$$3048 U$$3320/B1 U$$3054/A2 U$$719/B1 U$$3054/B2 VGND VGND VPWR VPWR U$$3049/A
+ sky130_fd_sc_hd__a22o_1
XU$$2314 _609_/Q U$$2318/A2 U$$2314/B1 U$$2318/B2 VGND VGND VPWR VPWR U$$2315/A sky130_fd_sc_hd__a22o_1
XU$$3059 U$$3059/A U$$3065/B VGND VGND VPWR VPWR U$$3059/X sky130_fd_sc_hd__xor2_1
XFILLER_46_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2325 U$$2325/A U$$2328/A VGND VGND VPWR VPWR U$$2325/X sky130_fd_sc_hd__xor2_1
XFILLER_62_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2336 U$$2336/A U$$2366/B VGND VGND VPWR VPWR U$$2336/X sky130_fd_sc_hd__xor2_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1602 U$$1602/A U$$1642/B VGND VGND VPWR VPWR U$$1602/X sky130_fd_sc_hd__xor2_1
XU$$2347 U$$429/A1 U$$2387/A2 U$$429/B1 U$$2387/B2 VGND VGND VPWR VPWR U$$2348/A sky130_fd_sc_hd__a22o_1
XU$$1613 U$$791/A1 U$$1627/A2 U$$517/B1 U$$1627/B2 VGND VGND VPWR VPWR U$$1614/A sky130_fd_sc_hd__a22o_1
XU$$2358 U$$2358/A U$$2388/B VGND VGND VPWR VPWR U$$2358/X sky130_fd_sc_hd__xor2_1
XU$$1624 U$$1624/A U$$1628/B VGND VGND VPWR VPWR U$$1624/X sky130_fd_sc_hd__xor2_1
XU$$2369 U$$2641/B1 U$$2423/A2 U$$2508/A1 U$$2423/B2 VGND VGND VPWR VPWR U$$2370/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1635 U$$950/A1 U$$1635/A2 U$$950/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1636/A sky130_fd_sc_hd__a22o_1
XU$$1646 _641_/Q VGND VGND VPWR VPWR U$$1646/Y sky130_fd_sc_hd__inv_1
XFILLER_188_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1657 U$$1657/A U$$1687/B VGND VGND VPWR VPWR U$$1657/X sky130_fd_sc_hd__xor2_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1668 U$$2077/B1 U$$1718/A2 U$$3312/B1 U$$1718/B2 VGND VGND VPWR VPWR U$$1669/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1679 U$$1679/A U$$1719/B VGND VGND VPWR VPWR U$$1679/X sky130_fd_sc_hd__xor2_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_308_ _444_/CLK _308_/D VGND VGND VPWR VPWR _308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_239_ _503_/CLK _239_/D VGND VGND VPWR VPWR _239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_61_2 dadda_fa_2_61_2/A dadda_fa_2_61_2/B dadda_fa_2_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/A dadda_fa_3_61_3/A sky130_fd_sc_hd__fa_1
Xrepeater502 U$$3066/A2 VGND VGND VPWR VPWR U$$3054/A2 sky130_fd_sc_hd__buf_4
XFILLER_57_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$309 final_adder.U$$308/A final_adder.U$$233/X final_adder.U$$235/X
+ VGND VGND VPWR VPWR final_adder.U$$309/X sky130_fd_sc_hd__a21o_1
Xrepeater513 U$$2981/A2 VGND VGND VPWR VPWR U$$2943/A2 sky130_fd_sc_hd__buf_6
Xrepeater524 U$$392/A2 VGND VGND VPWR VPWR U$$384/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_54_1 dadda_fa_2_54_1/A dadda_fa_2_54_1/B dadda_fa_2_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_0/CIN dadda_fa_3_54_2/CIN sky130_fd_sc_hd__fa_2
Xrepeater535 U$$2707/A2 VGND VGND VPWR VPWR U$$2697/A2 sky130_fd_sc_hd__buf_6
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater546 U$$2530/A2 VGND VGND VPWR VPWR U$$2524/A2 sky130_fd_sc_hd__buf_4
XFILLER_38_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater557 U$$2451/A2 VGND VGND VPWR VPWR U$$2437/A2 sky130_fd_sc_hd__buf_8
Xdadda_fa_5_31_0 dadda_fa_5_31_0/A dadda_fa_5_31_0/B dadda_fa_5_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_32_0/A dadda_fa_6_31_0/CIN sky130_fd_sc_hd__fa_2
Xrepeater568 U$$2059/X VGND VGND VPWR VPWR U$$2135/A2 sky130_fd_sc_hd__buf_4
XFILLER_168_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4250 U$$4350/B U$$4250/B VGND VGND VPWR VPWR U$$4250/X sky130_fd_sc_hd__and2_1
Xdadda_fa_2_47_0 U$$2761/X U$$2894/X U$$3027/X VGND VGND VPWR VPWR dadda_fa_3_48_0/B
+ dadda_fa_3_47_2/B sky130_fd_sc_hd__fa_1
Xrepeater579 U$$2038/A2 VGND VGND VPWR VPWR U$$2028/A2 sky130_fd_sc_hd__buf_6
XU$$4261 _555_/Q U$$4347/A2 _556_/Q U$$4347/B2 VGND VGND VPWR VPWR U$$4262/A sky130_fd_sc_hd__a22o_1
XFILLER_93_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4272 U$$4272/A U$$4298/B VGND VGND VPWR VPWR U$$4272/X sky130_fd_sc_hd__xor2_1
XFILLER_81_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4283 U$$4418/B1 U$$4327/A2 U$$4285/A1 U$$4319/B2 VGND VGND VPWR VPWR U$$4284/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4294 U$$4294/A U$$4296/B VGND VGND VPWR VPWR U$$4294/X sky130_fd_sc_hd__xor2_1
XU$$3560 U$$3560/A U$$3561/A VGND VGND VPWR VPWR U$$3560/X sky130_fd_sc_hd__xor2_1
XU$$3571 U$$3571/A U$$3613/B VGND VGND VPWR VPWR U$$3571/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3582 U$$4404/A1 U$$3628/A2 U$$4404/B1 U$$3628/B2 VGND VGND VPWR VPWR U$$3583/A
+ sky130_fd_sc_hd__a22o_1
XU$$3593 U$$3593/A U$$3637/B VGND VGND VPWR VPWR U$$3593/X sky130_fd_sc_hd__xor2_1
XFILLER_52_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2870 U$$3281/A1 U$$2874/A2 U$$3283/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2871/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_8_1 U$$627/B input245/X dadda_ha_4_8_0/SUM VGND VGND VPWR VPWR dadda_fa_6_9_0/B
+ dadda_fa_7_8_0/A sky130_fd_sc_hd__fa_1
XU$$2881 U$$2879/Y _658_/Q U$$2877/A U$$2880/X U$$2877/Y VGND VGND VPWR VPWR U$$2881/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_178_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2892 U$$2892/A U$$2944/B VGND VGND VPWR VPWR U$$2892/X sky130_fd_sc_hd__xor2_1
XFILLER_90_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_76_2 dadda_fa_4_76_2/A dadda_fa_4_76_2/B dadda_fa_4_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/CIN dadda_fa_5_76_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_161_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_69_1 dadda_fa_4_69_1/A dadda_fa_4_69_1/B dadda_fa_4_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/B dadda_fa_5_69_1/B sky130_fd_sc_hd__fa_1
XFILLER_88_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_332 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_46_0 dadda_fa_7_46_0/A dadda_fa_7_46_0/B dadda_fa_7_46_0/CIN VGND VGND
+ VPWR VPWR _471_/D _342_/D sky130_fd_sc_hd__fa_1
XFILLER_103_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$704 U$$704/A U$$726/B VGND VGND VPWR VPWR U$$704/X sky130_fd_sc_hd__xor2_1
XFILLER_56_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$715 U$$715/A1 U$$765/A2 U$$715/B1 U$$765/B2 VGND VGND VPWR VPWR U$$716/A sky130_fd_sc_hd__a22o_1
X_590_ _596_/CLK _590_/D VGND VGND VPWR VPWR _590_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$726 U$$726/A U$$726/B VGND VGND VPWR VPWR U$$726/X sky130_fd_sc_hd__xor2_1
XU$$737 U$$874/A1 U$$747/A2 U$$876/A1 U$$747/B2 VGND VGND VPWR VPWR U$$738/A sky130_fd_sc_hd__a22o_1
XFILLER_16_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$748 U$$748/A U$$748/B VGND VGND VPWR VPWR U$$748/X sky130_fd_sc_hd__xor2_1
XU$$759 U$$759/A1 U$$759/A2 U$$896/B1 U$$759/B2 VGND VGND VPWR VPWR U$$760/A sky130_fd_sc_hd__a22o_1
XFILLER_186_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1604 U$$32/A1 VGND VGND VPWR VPWR U$$991/A1 sky130_fd_sc_hd__buf_6
XANTENNA_9 ANTENNA_9/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1615 U$$3453/B1 VGND VGND VPWR VPWR U$$2494/B1 sky130_fd_sc_hd__buf_6
Xrepeater1626 _562_/Q VGND VGND VPWR VPWR U$$3042/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1637 U$$981/B1 VGND VGND VPWR VPWR U$$2077/B1 sky130_fd_sc_hd__buf_6
Xrepeater1648 U$$2625/A1 VGND VGND VPWR VPWR U$$22/A1 sky130_fd_sc_hd__buf_4
XFILLER_4_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1659 U$$4404/A1 VGND VGND VPWR VPWR U$$3717/B1 sky130_fd_sc_hd__buf_4
XFILLER_180_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_71_1 dadda_fa_3_71_1/A dadda_fa_3_71_1/B dadda_fa_3_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_0/CIN dadda_fa_4_71_2/A sky130_fd_sc_hd__fa_1
XFILLER_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_64_0 dadda_fa_3_64_0/A dadda_fa_3_64_0/B dadda_fa_3_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_0/B dadda_fa_4_64_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_750 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2100 U$$2100/A U$$2108/B VGND VGND VPWR VPWR U$$2100/X sky130_fd_sc_hd__xor2_1
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2111 U$$3618/A1 U$$2189/A2 _577_/Q U$$2189/B2 VGND VGND VPWR VPWR U$$2112/A sky130_fd_sc_hd__a22o_1
XFILLER_63_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_100_1 dadda_fa_4_100_1/A dadda_fa_4_100_1/B dadda_fa_4_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/B dadda_fa_5_100_1/B sky130_fd_sc_hd__fa_1
XU$$2122 U$$2122/A U$$2136/B VGND VGND VPWR VPWR U$$2122/X sky130_fd_sc_hd__xor2_1
XU$$2133 U$$624/B1 U$$2135/A2 U$$491/A1 U$$2135/B2 VGND VGND VPWR VPWR U$$2134/A sky130_fd_sc_hd__a22o_1
XU$$2144 U$$2144/A U$$2144/B VGND VGND VPWR VPWR U$$2144/X sky130_fd_sc_hd__xor2_1
XU$$1410 U$$449/B1 U$$1428/A2 U$$316/A1 U$$1428/B2 VGND VGND VPWR VPWR U$$1411/A sky130_fd_sc_hd__a22o_1
XU$$2155 U$$3386/B1 U$$2189/A2 U$$3388/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2156/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1421 U$$1421/A U$$1459/B VGND VGND VPWR VPWR U$$1421/X sky130_fd_sc_hd__xor2_1
XU$$2166 U$$2166/A U$$2170/B VGND VGND VPWR VPWR U$$2166/X sky130_fd_sc_hd__xor2_1
XU$$1432 U$$3213/A1 U$$1478/A2 U$$749/A1 U$$1478/B2 VGND VGND VPWR VPWR U$$1433/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2177 U$$3273/A1 U$$2185/A2 U$$2314/B1 U$$2185/B2 VGND VGND VPWR VPWR U$$2178/A
+ sky130_fd_sc_hd__a22o_1
XU$$1443 U$$1443/A U$$1443/B VGND VGND VPWR VPWR U$$1443/X sky130_fd_sc_hd__xor2_1
XU$$2188 U$$2188/A U$$2191/A VGND VGND VPWR VPWR U$$2188/X sky130_fd_sc_hd__xor2_1
XFILLER_16_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_499 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1454 U$$3096/B1 U$$1478/A2 U$$2415/A1 U$$1478/B2 VGND VGND VPWR VPWR U$$1455/A
+ sky130_fd_sc_hd__a22o_1
XU$$2199 U$$2199/A U$$2243/B VGND VGND VPWR VPWR U$$2199/X sky130_fd_sc_hd__xor2_1
XU$$1465 U$$1465/A U$$1475/B VGND VGND VPWR VPWR U$$1465/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1476 U$$2435/A1 U$$1374/X U$$791/B1 U$$1375/X VGND VGND VPWR VPWR U$$1477/A sky130_fd_sc_hd__a22o_1
XU$$1487 U$$1487/A U$$1487/B VGND VGND VPWR VPWR U$$1487/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_121_0 dadda_fa_7_121_0/A dadda_fa_7_121_0/B dadda_fa_7_121_0/CIN VGND
+ VGND VPWR VPWR _546_/D _417_/D sky130_fd_sc_hd__fa_1
XFILLER_31_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1498 U$$948/B1 U$$1500/A2 U$$952/A1 U$$1500/B2 VGND VGND VPWR VPWR U$$1499/A sky130_fd_sc_hd__a22o_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_86_1 dadda_fa_5_86_1/A dadda_fa_5_86_1/B dadda_fa_5_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_87_0/B dadda_fa_7_86_0/A sky130_fd_sc_hd__fa_2
XFILLER_144_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_79_0 dadda_fa_5_79_0/A dadda_fa_5_79_0/B dadda_fa_5_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_80_0/A dadda_fa_6_79_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_78_8 U$$4419/X input232/X dadda_fa_1_78_8/CIN VGND VGND VPWR VPWR dadda_fa_2_79_3/A
+ dadda_fa_3_78_0/A sky130_fd_sc_hd__fa_2
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$106 _530_/Q _402_/Q VGND VGND VPWR VPWR final_adder.U$$601/B1 final_adder.U$$728/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$117 _541_/Q _413_/Q VGND VGND VPWR VPWR final_adder.U$$245/B1 final_adder.U$$739/A
+ sky130_fd_sc_hd__ha_2
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$139 final_adder.U$$633/A final_adder.U$$505/B1 final_adder.U$$139/B1
+ VGND VGND VPWR VPWR final_adder.U$$139/X sky130_fd_sc_hd__a21o_1
Xrepeater387 U$$999/A2 VGND VGND VPWR VPWR U$$1039/A2 sky130_fd_sc_hd__buf_4
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater398 U$$948/A2 VGND VGND VPWR VPWR U$$924/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4080 U$$4080/A U$$4084/B VGND VGND VPWR VPWR U$$4080/X sky130_fd_sc_hd__xor2_1
XFILLER_66_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4091 U$$4500/B1 U$$4095/A2 U$$4228/B1 U$$4105/B2 VGND VGND VPWR VPWR U$$4092/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3390 _599_/Q U$$3402/A2 _600_/Q U$$3402/B2 VGND VGND VPWR VPWR U$$3391/A sky130_fd_sc_hd__a22o_1
XFILLER_0_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_81_0 dadda_fa_4_81_0/A dadda_fa_4_81_0/B dadda_fa_4_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/A dadda_fa_5_81_1/A sky130_fd_sc_hd__fa_1
XFILLER_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_102_3 dadda_fa_3_102_3/A dadda_fa_3_102_3/B dadda_fa_3_102_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_103_1/B dadda_fa_4_102_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput102 b[43] VGND VGND VPWR VPWR _595_/D sky130_fd_sc_hd__clkbuf_1
Xinput113 b[53] VGND VGND VPWR VPWR _605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput124 b[63] VGND VGND VPWR VPWR _615_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput135 c[105] VGND VGND VPWR VPWR input135/X sky130_fd_sc_hd__buf_2
XTAP_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput146 c[115] VGND VGND VPWR VPWR input146/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput157 c[125] VGND VGND VPWR VPWR input157/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 c[1] VGND VGND VPWR VPWR input168/X sky130_fd_sc_hd__clkbuf_4
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 c[2] VGND VGND VPWR VPWR input179/X sky130_fd_sc_hd__clkbuf_4
Xfinal_adder.U$$640 final_adder.U$$640/A final_adder.U$$640/B VGND VGND VPWR VPWR
+ _186_/D sky130_fd_sc_hd__xor2_4
XTAP_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_642_ _642_/CLK _642_/D VGND VGND VPWR VPWR _642_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$651 final_adder.U$$651/A final_adder.U$$651/B VGND VGND VPWR VPWR
+ _197_/D sky130_fd_sc_hd__xor2_4
XFILLER_91_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$662 final_adder.U$$662/A final_adder.U$$662/B VGND VGND VPWR VPWR
+ _208_/D sky130_fd_sc_hd__xor2_1
XTAP_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_109_0 dadda_fa_6_109_0/A dadda_fa_6_109_0/B dadda_fa_6_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_110_0/B dadda_fa_7_109_0/CIN sky130_fd_sc_hd__fa_1
XU$$501 U$$501/A1 U$$517/A2 U$$912/B1 U$$517/B2 VGND VGND VPWR VPWR U$$502/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$673 final_adder.U$$673/A final_adder.U$$673/B VGND VGND VPWR VPWR
+ _219_/D sky130_fd_sc_hd__xor2_1
XTAP_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$512 U$$512/A U$$518/B VGND VGND VPWR VPWR U$$512/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$684 final_adder.U$$684/A final_adder.U$$684/B VGND VGND VPWR VPWR
+ _230_/D sky130_fd_sc_hd__xor2_1
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$523 U$$658/B1 U$$545/A2 U$$525/A1 U$$545/B2 VGND VGND VPWR VPWR U$$524/A sky130_fd_sc_hd__a22o_1
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$695 final_adder.U$$695/A final_adder.U$$695/B VGND VGND VPWR VPWR
+ _241_/D sky130_fd_sc_hd__xor2_2
XU$$534 U$$534/A U$$536/B VGND VGND VPWR VPWR U$$534/X sky130_fd_sc_hd__xor2_1
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_573_ _575_/CLK _573_/D VGND VGND VPWR VPWR _573_/Q sky130_fd_sc_hd__dfxtp_4
XU$$545 U$$545/A1 U$$545/A2 U$$545/B1 U$$545/B2 VGND VGND VPWR VPWR U$$546/A sky130_fd_sc_hd__a22o_1
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$556 U$$828/B1 U$$600/A2 U$$556/B1 U$$600/B2 VGND VGND VPWR VPWR U$$557/A sky130_fd_sc_hd__a22o_1
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$567 U$$567/A U$$589/B VGND VGND VPWR VPWR U$$567/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_29_3 dadda_fa_3_29_3/A dadda_fa_3_29_3/B dadda_fa_3_29_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_30_1/B dadda_fa_4_29_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_44_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$578 U$$715/A1 U$$600/A2 U$$715/B1 U$$600/B2 VGND VGND VPWR VPWR U$$579/A sky130_fd_sc_hd__a22o_1
XU$$589 U$$589/A U$$589/B VGND VGND VPWR VPWR U$$589/X sky130_fd_sc_hd__xor2_1
XFILLER_189_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_96_0 dadda_fa_6_96_0/A dadda_fa_6_96_0/B dadda_fa_6_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_97_0/B dadda_fa_7_96_0/CIN sky130_fd_sc_hd__fa_1
Xclkbuf_3_1__f_clk clkbuf_2_0_0_clk/X VGND VGND VPWR VPWR _616_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_201_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1401 U$$4468/A1 VGND VGND VPWR VPWR U$$3646/A1 sky130_fd_sc_hd__buf_6
XFILLER_193_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1412 U$$4053/A1 VGND VGND VPWR VPWR U$$900/B1 sky130_fd_sc_hd__buf_4
Xrepeater1423 _587_/Q VGND VGND VPWR VPWR U$$4051/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1434 _586_/Q VGND VGND VPWR VPWR U$$4323/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1445 U$$4317/B1 VGND VGND VPWR VPWR U$$2947/B1 sky130_fd_sc_hd__buf_6
XFILLER_67_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1456 U$$3769/A1 VGND VGND VPWR VPWR U$$890/B1 sky130_fd_sc_hd__buf_4
XFILLER_180_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1467 U$$4450/A1 VGND VGND VPWR VPWR U$$3217/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_153_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1478 U$$4448/A1 VGND VGND VPWR VPWR U$$201/A1 sky130_fd_sc_hd__buf_6
XFILLER_119_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1489 U$$4444/B1 VGND VGND VPWR VPWR U$$4035/A1 sky130_fd_sc_hd__buf_4
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_2_32_5 U$$2066/X U$$2199/X VGND VGND VPWR VPWR dadda_fa_3_33_2/A dadda_fa_4_32_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_80_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_31_3 U$$1266/X U$$1399/X U$$1532/X VGND VGND VPWR VPWR dadda_fa_3_32_1/CIN
+ dadda_fa_3_31_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_208_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1240 U$$1240/A U$$1288/B VGND VGND VPWR VPWR U$$1240/X sky130_fd_sc_hd__xor2_1
XU$$1251 U$$429/A1 U$$1295/A2 U$$429/B1 U$$1295/B2 VGND VGND VPWR VPWR U$$1252/A sky130_fd_sc_hd__a22o_1
XU$$1262 U$$1262/A U$$1292/B VGND VGND VPWR VPWR U$$1262/X sky130_fd_sc_hd__xor2_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1273 U$$2641/B1 U$$1279/A2 U$$2508/A1 U$$1279/B2 VGND VGND VPWR VPWR U$$1274/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1284 U$$1284/A U$$1292/B VGND VGND VPWR VPWR U$$1284/X sky130_fd_sc_hd__xor2_1
XFILLER_31_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1295 U$$3213/A1 U$$1295/A2 U$$749/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1296/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_83_6 U$$3764/X U$$3897/X U$$4030/X VGND VGND VPWR VPWR dadda_fa_2_84_3/CIN
+ dadda_fa_3_83_0/A sky130_fd_sc_hd__fa_1
XFILLER_171_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_76_5 U$$3484/X U$$3617/X U$$3750/X VGND VGND VPWR VPWR dadda_fa_2_77_2/A
+ dadda_fa_2_76_5/A sky130_fd_sc_hd__fa_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_4 U$$4002/X U$$4135/X U$$4268/X VGND VGND VPWR VPWR dadda_fa_2_70_1/CIN
+ dadda_fa_2_69_4/CIN sky130_fd_sc_hd__fa_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_39_2 dadda_fa_4_39_2/A dadda_fa_4_39_2/B dadda_fa_4_39_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/CIN dadda_fa_5_39_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_207 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_229 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_100_0 U$$4330/X U$$4463/X input130/X VGND VGND VPWR VPWR dadda_fa_4_101_0/B
+ dadda_fa_4_100_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_64_3 U$$1332/X U$$1465/X U$$1598/X VGND VGND VPWR VPWR dadda_fa_1_65_6/B
+ dadda_fa_1_64_8/B sky130_fd_sc_hd__fa_1
XFILLER_77_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$0_1711 VGND VGND VPWR VPWR U$$0_1711/HI U$$0/A sky130_fd_sc_hd__conb_1
Xdadda_fa_3_41_2 dadda_fa_3_41_2/A dadda_fa_3_41_2/B dadda_fa_3_41_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_1/A dadda_fa_4_41_2/B sky130_fd_sc_hd__fa_2
XTAP_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$481 final_adder.U$$304/B final_adder.U$$718/B final_adder.U$$225/X
+ VGND VGND VPWR VPWR final_adder.U$$720/B sky130_fd_sc_hd__a21o_1
XFILLER_205_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_34_1 dadda_fa_3_34_1/A dadda_fa_3_34_1/B dadda_fa_3_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_0/CIN dadda_fa_4_34_2/A sky130_fd_sc_hd__fa_1
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_625_ _633_/CLK _625_/D VGND VGND VPWR VPWR _625_/Q sky130_fd_sc_hd__dfxtp_1
XU$$320 U$$729/B1 U$$334/A2 U$$733/A1 U$$334/B2 VGND VGND VPWR VPWR U$$321/A sky130_fd_sc_hd__a22o_1
XFILLER_91_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$331 U$$331/A U$$397/B VGND VGND VPWR VPWR U$$331/X sky130_fd_sc_hd__xor2_1
XU$$342 U$$614/B1 U$$350/A2 U$$344/A1 U$$350/B2 VGND VGND VPWR VPWR U$$343/A sky130_fd_sc_hd__a22o_1
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$353 U$$353/A U$$397/B VGND VGND VPWR VPWR U$$353/X sky130_fd_sc_hd__xor2_1
XFILLER_33_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_11_0 dadda_fa_6_11_0/A dadda_fa_6_11_0/B dadda_fa_6_11_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_12_0/B dadda_fa_7_11_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_27_0 U$$1125/X U$$1258/X U$$1391/X VGND VGND VPWR VPWR dadda_fa_4_28_0/B
+ dadda_fa_4_27_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_33_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_926 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$364 U$$501/A1 U$$392/A2 U$$912/B1 U$$392/B2 VGND VGND VPWR VPWR U$$365/A sky130_fd_sc_hd__a22o_1
XFILLER_205_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$375 U$$375/A U$$383/B VGND VGND VPWR VPWR U$$375/X sky130_fd_sc_hd__xor2_1
X_556_ _558_/CLK _556_/D VGND VGND VPWR VPWR _556_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$386 U$$658/B1 U$$392/A2 U$$525/A1 U$$392/B2 VGND VGND VPWR VPWR U$$387/A sky130_fd_sc_hd__a22o_1
XU$$397 U$$397/A U$$397/B VGND VGND VPWR VPWR U$$397/X sky130_fd_sc_hd__xor2_1
XFILLER_33_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_487_ _487_/CLK _487_/D VGND VGND VPWR VPWR _487_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_186_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_93_5 dadda_fa_2_93_5/A dadda_fa_2_93_5/B dadda_fa_2_93_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_94_2/A dadda_fa_4_93_0/A sky130_fd_sc_hd__fa_2
Xrepeater1220 U$$3551/B1 VGND VGND VPWR VPWR U$$4512/A1 sky130_fd_sc_hd__buf_4
Xrepeater1231 _611_/Q VGND VGND VPWR VPWR U$$2866/A1 sky130_fd_sc_hd__buf_6
XFILLER_99_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1242 U$$2725/A1 VGND VGND VPWR VPWR U$$2586/B1 sky130_fd_sc_hd__buf_6
Xrepeater1253 U$$3269/B1 VGND VGND VPWR VPWR U$$940/B1 sky130_fd_sc_hd__buf_6
Xrepeater1264 _607_/Q VGND VGND VPWR VPWR U$$3132/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_86_4 dadda_fa_2_86_4/A dadda_fa_2_86_4/B dadda_fa_2_86_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_1/CIN dadda_fa_3_86_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1275 U$$2717/A1 VGND VGND VPWR VPWR U$$525/A1 sky130_fd_sc_hd__clkbuf_8
Xrepeater1286 U$$4222/A1 VGND VGND VPWR VPWR U$$4494/B1 sky130_fd_sc_hd__buf_6
XFILLER_180_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1297 _603_/Q VGND VGND VPWR VPWR U$$3807/B1 sky130_fd_sc_hd__buf_4
XFILLER_114_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_79_3 dadda_fa_2_79_3/A dadda_fa_2_79_3/B dadda_fa_2_79_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/B dadda_fa_3_79_3/B sky130_fd_sc_hd__fa_1
XFILLER_45_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1367_1717 VGND VGND VPWR VPWR U$$1367_1717/HI U$$1367/B1 sky130_fd_sc_hd__conb_1
XFILLER_171_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_49_1 dadda_fa_5_49_1/A dadda_fa_5_49_1/B dadda_fa_5_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_50_0/B dadda_fa_7_49_0/A sky130_fd_sc_hd__fa_1
XFILLER_110_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_336 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_102_2 U$$3403/X U$$3536/X U$$3669/X VGND VGND VPWR VPWR dadda_fa_3_103_2/CIN
+ dadda_fa_3_102_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_51_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1070 U$$1070/A _631_/Q VGND VGND VPWR VPWR U$$1070/X sky130_fd_sc_hd__xor2_1
XFILLER_143_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1081 U$$942/B1 U$$1093/A2 U$$2588/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1082/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1092 U$$1092/A U$$1095/A VGND VGND VPWR VPWR U$$1092/X sky130_fd_sc_hd__xor2_1
XFILLER_32_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_806 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_123_1 U$$4509/X input155/X dadda_fa_5_123_1/CIN VGND VGND VPWR VPWR dadda_fa_6_124_0/B
+ dadda_fa_7_123_0/A sky130_fd_sc_hd__fa_1
XFILLER_31_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2326_1732 VGND VGND VPWR VPWR U$$2326_1732/HI U$$2326/B1 sky130_fd_sc_hd__conb_1
Xdadda_fa_5_116_0 dadda_fa_5_116_0/A dadda_fa_5_116_0/B dadda_fa_5_116_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_117_0/A dadda_fa_6_116_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_81_3 U$$2430/X U$$2563/X U$$2696/X VGND VGND VPWR VPWR dadda_fa_2_82_2/A
+ dadda_fa_2_81_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_137_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_74_2 U$$2549/X U$$2682/X U$$2815/X VGND VGND VPWR VPWR dadda_fa_2_75_1/A
+ dadda_fa_2_74_4/A sky130_fd_sc_hd__fa_1
XFILLER_137_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_51_1 dadda_fa_4_51_1/A dadda_fa_4_51_1/B dadda_fa_4_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/B dadda_fa_5_51_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_67_1 U$$2934/X U$$3067/X U$$3200/X VGND VGND VPWR VPWR dadda_fa_2_68_0/CIN
+ dadda_fa_2_67_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_44_0 dadda_fa_4_44_0/A dadda_fa_4_44_0/B dadda_fa_4_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/A dadda_fa_5_44_1/A sky130_fd_sc_hd__fa_1
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1067 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_410_ _648_/CLK _410_/D VGND VGND VPWR VPWR _410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_341_ _470_/CLK _341_/D VGND VGND VPWR VPWR _341_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_272_ _521_/CLK _272_/D VGND VGND VPWR VPWR _272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_96_3 dadda_fa_3_96_3/A dadda_fa_3_96_3/B dadda_fa_3_96_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_1/B dadda_fa_4_96_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_6_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_89_2 dadda_fa_3_89_2/A dadda_fa_3_89_2/B dadda_fa_3_89_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_1/A dadda_fa_4_89_2/B sky130_fd_sc_hd__fa_1
XFILLER_159_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_59_0 dadda_fa_6_59_0/A dadda_fa_6_59_0/B dadda_fa_6_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_60_0/B dadda_fa_7_59_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_78_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater909 _679_/Q VGND VGND VPWR VPWR U$$4350/B sky130_fd_sc_hd__buf_6
Xdadda_fa_0_62_0 U$$131/X U$$264/X U$$397/X VGND VGND VPWR VPWR dadda_fa_1_63_5/B
+ dadda_fa_1_62_7/B sky130_fd_sc_hd__fa_2
XFILLER_65_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3901 U$$3901/A U$$3949/B VGND VGND VPWR VPWR U$$3901/X sky130_fd_sc_hd__xor2_1
XFILLER_77_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3912 U$$4323/A1 U$$3932/A2 U$$4462/A1 U$$3932/B2 VGND VGND VPWR VPWR U$$3913/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3923 U$$3923/A U$$3935/B VGND VGND VPWR VPWR U$$3923/X sky130_fd_sc_hd__xor2_1
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3934 U$$4206/B1 U$$3840/X U$$3934/B1 U$$3841/X VGND VGND VPWR VPWR U$$3935/A sky130_fd_sc_hd__a22o_1
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3945 U$$3945/A U$$3949/B VGND VGND VPWR VPWR U$$3945/X sky130_fd_sc_hd__xor2_1
XU$$3956 U$$4228/B1 U$$3958/A2 U$$4369/A1 U$$3958/B2 VGND VGND VPWR VPWR U$$3957/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3967 U$$3967/A U$$3973/A VGND VGND VPWR VPWR U$$3967/X sky130_fd_sc_hd__xor2_1
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3978 U$$3976/B _673_/Q _674_/Q U$$3973/Y VGND VGND VPWR VPWR U$$3978/X sky130_fd_sc_hd__a22o_1
X_608_ _613_/CLK _608_/D VGND VGND VPWR VPWR _608_/Q sky130_fd_sc_hd__dfxtp_2
XU$$150 U$$150/A U$$180/B VGND VGND VPWR VPWR U$$150/X sky130_fd_sc_hd__xor2_1
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3989 U$$4400/A1 U$$4005/A2 U$$4402/A1 U$$4005/B2 VGND VGND VPWR VPWR U$$3990/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$161 U$$22/B1 U$$175/A2 U$$26/A1 U$$175/B2 VGND VGND VPWR VPWR U$$162/A sky130_fd_sc_hd__a22o_1
XU$$172 U$$172/A U$$196/B VGND VGND VPWR VPWR U$$172/X sky130_fd_sc_hd__xor2_1
XFILLER_72_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$183 U$$866/B1 U$$219/A2 U$$733/A1 U$$219/B2 VGND VGND VPWR VPWR U$$184/A sky130_fd_sc_hd__a22o_1
XU$$194 U$$194/A U$$196/B VGND VGND VPWR VPWR U$$194/X sky130_fd_sc_hd__xor2_1
XFILLER_36_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_539_ _648_/CLK _539_/D VGND VGND VPWR VPWR _539_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_496 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_91_2 U$$3913/X U$$4046/X U$$4179/X VGND VGND VPWR VPWR dadda_fa_3_92_1/A
+ dadda_fa_3_91_3/A sky130_fd_sc_hd__fa_1
XFILLER_126_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1050 U$$2144/B VGND VGND VPWR VPWR U$$2110/B sky130_fd_sc_hd__buf_6
Xrepeater1061 U$$2043/B VGND VGND VPWR VPWR U$$2039/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_84_1 U$$4431/X input239/X dadda_fa_2_84_1/CIN VGND VGND VPWR VPWR dadda_fa_3_85_0/CIN
+ dadda_fa_3_84_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput258 _268_/Q VGND VGND VPWR VPWR o[100] sky130_fd_sc_hd__buf_2
Xrepeater1072 U$$1918/A VGND VGND VPWR VPWR U$$1916/B sky130_fd_sc_hd__buf_6
XFILLER_86_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1083 U$$1554/B VGND VGND VPWR VPWR U$$1558/B sky130_fd_sc_hd__buf_8
Xoutput269 _278_/Q VGND VGND VPWR VPWR o[110] sky130_fd_sc_hd__buf_2
Xdadda_fa_5_61_0 dadda_fa_5_61_0/A dadda_fa_5_61_0/B dadda_fa_5_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_62_0/A dadda_fa_6_61_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1094 _637_/Q VGND VGND VPWR VPWR U$$1475/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_77_0 dadda_fa_2_77_0/A dadda_fa_2_77_0/B dadda_fa_2_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_0/B dadda_fa_3_77_2/B sky130_fd_sc_hd__fa_1
XFILLER_142_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1230_1714 VGND VGND VPWR VPWR U$$1230_1714/HI U$$1230/B1 sky130_fd_sc_hd__conb_1
XFILLER_99_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_60_8 dadda_fa_1_60_8/A dadda_fa_1_60_8/B dadda_fa_1_60_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_61_3/A dadda_fa_3_60_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_1_53_7 U$$3172/X U$$3305/X U$$3438/X VGND VGND VPWR VPWR dadda_fa_2_54_2/CIN
+ dadda_fa_2_53_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_56_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4443_1800 VGND VGND VPWR VPWR U$$4443_1800/HI U$$4443/B sky130_fd_sc_hd__conb_1
XFILLER_208_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1023 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_444 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_99_1 dadda_fa_4_99_1/A dadda_fa_4_99_1/B dadda_fa_4_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/B dadda_fa_5_99_1/B sky130_fd_sc_hd__fa_1
XFILLER_152_606 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_76_0 dadda_fa_7_76_0/A dadda_fa_7_76_0/B dadda_fa_7_76_0/CIN VGND VGND
+ VPWR VPWR _501_/D _372_/D sky130_fd_sc_hd__fa_1
XFILLER_191_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_371 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3208 U$$3208/A U$$3208/B VGND VGND VPWR VPWR U$$3208/X sky130_fd_sc_hd__xor2_1
XU$$3219 U$$3354/B1 U$$3263/A2 U$$3221/A1 U$$3263/B2 VGND VGND VPWR VPWR U$$3220/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1038 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2507 U$$2507/A U$$2551/B VGND VGND VPWR VPWR U$$2507/X sky130_fd_sc_hd__xor2_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2518 U$$3475/B1 U$$2524/A2 U$$3342/A1 U$$2524/B2 VGND VGND VPWR VPWR U$$2519/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2529 U$$2529/A U$$2531/B VGND VGND VPWR VPWR U$$2529/X sky130_fd_sc_hd__xor2_1
XFILLER_62_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1806 U$$1806/A U$$1844/B VGND VGND VPWR VPWR U$$1806/X sky130_fd_sc_hd__xor2_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1817 U$$36/A1 U$$1859/A2 U$$38/A1 U$$1859/B2 VGND VGND VPWR VPWR U$$1818/A sky130_fd_sc_hd__a22o_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1828 U$$1828/A U$$1874/B VGND VGND VPWR VPWR U$$1828/X sky130_fd_sc_hd__xor2_1
XU$$1839 U$$1976/A1 U$$1843/A2 U$$3485/A1 U$$1843/B2 VGND VGND VPWR VPWR U$$1840/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_324_ _469_/CLK _324_/D VGND VGND VPWR VPWR _324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_255_ _379_/CLK _255_/D VGND VGND VPWR VPWR _255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_186_ _189_/CLK _186_/D VGND VGND VPWR VPWR _186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_94_0 dadda_fa_3_94_0/A dadda_fa_3_94_0/B dadda_fa_3_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_0/B dadda_fa_4_94_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4390_1773 VGND VGND VPWR VPWR U$$4390_1773/HI U$$4390/A1 sky130_fd_sc_hd__conb_1
XFILLER_69_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater706 U$$3841/X VGND VGND VPWR VPWR U$$3910/B2 sky130_fd_sc_hd__buf_6
XFILLER_42_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater717 U$$3704/X VGND VGND VPWR VPWR U$$3805/B2 sky130_fd_sc_hd__buf_6
Xrepeater728 U$$3537/B2 VGND VGND VPWR VPWR U$$3519/B2 sky130_fd_sc_hd__buf_4
XU$$4410 U$$4410/A1 U$$4388/X _562_/Q U$$4430/B2 VGND VGND VPWR VPWR U$$4411/A sky130_fd_sc_hd__a22o_1
XFILLER_42_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_56_5 dadda_fa_2_56_5/A dadda_fa_2_56_5/B dadda_fa_2_56_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_2/A dadda_fa_4_56_0/A sky130_fd_sc_hd__fa_2
XU$$4421 U$$4421/A U$$4421/B VGND VGND VPWR VPWR U$$4421/X sky130_fd_sc_hd__xor2_1
XFILLER_65_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater739 U$$3404/B2 VGND VGND VPWR VPWR U$$3402/B2 sky130_fd_sc_hd__buf_6
XU$$4432 U$$4432/A1 U$$4388/X U$$4434/A1 U$$4438/B2 VGND VGND VPWR VPWR U$$4433/A
+ sky130_fd_sc_hd__a22o_1
XU$$4443 U$$4443/A U$$4443/B VGND VGND VPWR VPWR U$$4443/X sky130_fd_sc_hd__xor2_1
XU$$4454 _583_/Q U$$4388/X _584_/Q U$$4454/B2 VGND VGND VPWR VPWR U$$4455/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_4 dadda_fa_2_49_4/A dadda_fa_2_49_4/B dadda_fa_2_49_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/CIN dadda_fa_3_49_3/CIN sky130_fd_sc_hd__fa_1
XU$$4465 U$$4465/A U$$4465/B VGND VGND VPWR VPWR U$$4465/X sky130_fd_sc_hd__xor2_1
XU$$3720 U$$3720/A U$$3740/B VGND VGND VPWR VPWR U$$3720/X sky130_fd_sc_hd__xor2_1
XFILLER_93_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3731 _564_/Q U$$3769/A2 _565_/Q U$$3769/B2 VGND VGND VPWR VPWR U$$3732/A sky130_fd_sc_hd__a22o_1
XU$$4476 U$$4476/A1 U$$4388/X U$$4478/A1 U$$4480/B2 VGND VGND VPWR VPWR U$$4477/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4487 U$$4487/A U$$4487/B VGND VGND VPWR VPWR U$$4487/X sky130_fd_sc_hd__xor2_1
XU$$3742 U$$3742/A U$$3764/B VGND VGND VPWR VPWR U$$3742/X sky130_fd_sc_hd__xor2_1
XU$$3753 U$$3753/A1 U$$3785/A2 _576_/Q U$$3785/B2 VGND VGND VPWR VPWR U$$3754/A sky130_fd_sc_hd__a22o_1
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4498 U$$4498/A1 U$$4388/X U$$938/A1 U$$4389/X VGND VGND VPWR VPWR U$$4499/A sky130_fd_sc_hd__a22o_1
XFILLER_65_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3764 U$$3764/A U$$3764/B VGND VGND VPWR VPWR U$$3764/X sky130_fd_sc_hd__xor2_1
XU$$3775 U$$4323/A1 U$$3777/A2 U$$4462/A1 U$$3777/B2 VGND VGND VPWR VPWR U$$3776/A
+ sky130_fd_sc_hd__a22o_1
XU$$3786 U$$3786/A U$$3800/B VGND VGND VPWR VPWR U$$3786/X sky130_fd_sc_hd__xor2_1
XFILLER_46_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3797 U$$4206/B1 U$$3805/A2 U$$3934/B1 U$$3805/B2 VGND VGND VPWR VPWR U$$3798/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_390 _569_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$622_1848 VGND VGND VPWR VPWR final_adder.U$$622_1848/HI final_adder.U$$622/B
+ sky130_fd_sc_hd__conb_1
XFILLER_119_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_934 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4473_1815 VGND VGND VPWR VPWR U$$4473_1815/HI U$$4473/B sky130_fd_sc_hd__conb_1
XFILLER_109_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_45_5 U$$2092/X U$$2225/X VGND VGND VPWR VPWR dadda_fa_2_46_3/CIN dadda_fa_3_45_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_87_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_51_4 U$$1705/X U$$1838/X U$$1971/X VGND VGND VPWR VPWR dadda_fa_2_52_1/CIN
+ dadda_fa_2_51_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$908 U$$908/A1 U$$956/A2 U$$910/A1 U$$956/B2 VGND VGND VPWR VPWR U$$909/A sky130_fd_sc_hd__a22o_1
XU$$919 U$$919/A U$$951/B VGND VGND VPWR VPWR U$$919/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_44_3 U$$1292/X U$$1425/X U$$1558/X VGND VGND VPWR VPWR dadda_fa_2_45_3/B
+ dadda_fa_2_44_5/B sky130_fd_sc_hd__fa_1
XFILLER_44_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_21_2 dadda_fa_4_21_2/A dadda_fa_4_21_2/B dadda_ha_3_21_3/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_22_0/CIN dadda_fa_5_21_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_14_1 U$$700/X U$$833/X U$$966/X VGND VGND VPWR VPWR dadda_fa_5_15_0/B
+ dadda_fa_5_14_1/B sky130_fd_sc_hd__fa_1
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1014 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_5_126_0_1878 VGND VGND VPWR VPWR dadda_ha_5_126_0/A dadda_ha_5_126_0_1878/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_59_3 dadda_fa_3_59_3/A dadda_fa_3_59_3/B dadda_fa_3_59_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_1/B dadda_fa_4_59_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3005 U$$3005/A1 U$$3005/A2 U$$3281/A1 U$$3005/B2 VGND VGND VPWR VPWR U$$3006/A
+ sky130_fd_sc_hd__a22o_1
XU$$3016 _661_/Q VGND VGND VPWR VPWR U$$3016/Y sky130_fd_sc_hd__inv_1
XFILLER_208_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3027 U$$3027/A U$$3077/B VGND VGND VPWR VPWR U$$3027/X sky130_fd_sc_hd__xor2_1
XU$$3038 U$$3175/A1 U$$3046/A2 U$$4410/A1 U$$3046/B2 VGND VGND VPWR VPWR U$$3039/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2304 U$$4494/B1 U$$2196/X U$$4224/A1 U$$2197/X VGND VGND VPWR VPWR U$$2305/A sky130_fd_sc_hd__a22o_1
XFILLER_74_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3049 U$$3049/A U$$3049/B VGND VGND VPWR VPWR U$$3049/X sky130_fd_sc_hd__xor2_1
XU$$2315 U$$2315/A U$$2321/B VGND VGND VPWR VPWR U$$2315/X sky130_fd_sc_hd__xor2_1
XU$$2326 U$$956/A1 U$$2326/A2 U$$2326/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2327/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2337 U$$2611/A1 U$$2367/A2 U$$2611/B1 U$$2367/B2 VGND VGND VPWR VPWR U$$2338/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1603 U$$2971/B1 U$$1607/A2 U$$2838/A1 U$$1607/B2 VGND VGND VPWR VPWR U$$1604/A
+ sky130_fd_sc_hd__a22o_1
XU$$2348 U$$2348/A U$$2388/B VGND VGND VPWR VPWR U$$2348/X sky130_fd_sc_hd__xor2_1
XFILLER_90_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1614 U$$1614/A U$$1628/B VGND VGND VPWR VPWR U$$1614/X sky130_fd_sc_hd__xor2_1
XFILLER_188_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2359 U$$2494/B1 U$$2387/A2 U$$854/A1 U$$2387/B2 VGND VGND VPWR VPWR U$$2360/A
+ sky130_fd_sc_hd__a22o_1
XU$$1625 U$$2858/A1 U$$1627/A2 U$$2721/B1 U$$1627/B2 VGND VGND VPWR VPWR U$$1626/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1636 U$$1636/A U$$1636/B VGND VGND VPWR VPWR U$$1636/X sky130_fd_sc_hd__xor2_1
XU$$1647 _641_/Q U$$1647/B VGND VGND VPWR VPWR U$$1647/X sky130_fd_sc_hd__and2_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1658 U$$973/A1 U$$1684/A2 U$$838/A1 U$$1684/B2 VGND VGND VPWR VPWR U$$1659/A sky130_fd_sc_hd__a22o_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1669 U$$1669/A U$$1719/B VGND VGND VPWR VPWR U$$1669/X sky130_fd_sc_hd__xor2_1
XFILLER_15_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_307_ _435_/CLK _307_/D VGND VGND VPWR VPWR _307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_238_ _503_/CLK _238_/D VGND VGND VPWR VPWR _238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_169_ _179_/CLK _169_/D VGND VGND VPWR VPWR _169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_61_3 dadda_fa_2_61_3/A dadda_fa_2_61_3/B dadda_fa_2_61_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/B dadda_fa_3_61_3/B sky130_fd_sc_hd__fa_1
Xrepeater503 U$$3148/A2 VGND VGND VPWR VPWR U$$3066/A2 sky130_fd_sc_hd__buf_4
XFILLER_85_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater514 U$$3005/A2 VGND VGND VPWR VPWR U$$2959/A2 sky130_fd_sc_hd__buf_6
XFILLER_38_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater525 U$$408/A2 VGND VGND VPWR VPWR U$$392/A2 sky130_fd_sc_hd__buf_6
XFILLER_66_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_54_2 dadda_fa_2_54_2/A dadda_fa_2_54_2/B dadda_fa_2_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/A dadda_fa_3_54_3/A sky130_fd_sc_hd__fa_1
Xrepeater536 U$$2663/A2 VGND VGND VPWR VPWR U$$2653/A2 sky130_fd_sc_hd__buf_4
Xrepeater547 U$$2470/X VGND VGND VPWR VPWR U$$2530/A2 sky130_fd_sc_hd__buf_4
XU$$4240 U$$4514/A1 U$$4244/A2 U$$4516/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4241/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater558 U$$2333/X VGND VGND VPWR VPWR U$$2451/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_5_31_1 dadda_fa_5_31_1/A dadda_fa_5_31_1/B dadda_fa_5_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_32_0/B dadda_fa_7_31_0/A sky130_fd_sc_hd__fa_1
XU$$4251 U$$4249/Y _678_/Q U$$4247/A U$$4250/X U$$4247/Y VGND VGND VPWR VPWR U$$4251/X
+ sky130_fd_sc_hd__a32o_4
Xrepeater569 U$$2115/A2 VGND VGND VPWR VPWR U$$2109/A2 sky130_fd_sc_hd__buf_6
XFILLER_168_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4262 U$$4262/A U$$4384/A VGND VGND VPWR VPWR U$$4262/X sky130_fd_sc_hd__xor2_1
XFILLER_66_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_47_1 U$$3160/X input198/X dadda_fa_2_47_1/CIN VGND VGND VPWR VPWR dadda_fa_3_48_0/CIN
+ dadda_fa_3_47_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_26_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3559_1752 VGND VGND VPWR VPWR U$$3559_1752/HI U$$3559/B1 sky130_fd_sc_hd__conb_1
XU$$4273 U$$4273/A1 U$$4297/A2 U$$4273/B1 U$$4297/B2 VGND VGND VPWR VPWR U$$4274/A
+ sky130_fd_sc_hd__a22o_1
XU$$4284 U$$4284/A U$$4322/B VGND VGND VPWR VPWR U$$4284/X sky130_fd_sc_hd__xor2_1
XFILLER_81_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_24_0 dadda_fa_5_24_0/A dadda_fa_5_24_0/B dadda_fa_5_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_25_0/A dadda_fa_6_24_0/CIN sky130_fd_sc_hd__fa_1
XU$$3550 U$$3550/A U$$3556/B VGND VGND VPWR VPWR U$$3550/X sky130_fd_sc_hd__xor2_1
XFILLER_52_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4295 U$$4432/A1 U$$4311/A2 _573_/Q U$$4311/B2 VGND VGND VPWR VPWR U$$4296/A sky130_fd_sc_hd__a22o_1
XU$$3561 U$$3561/A VGND VGND VPWR VPWR U$$3561/Y sky130_fd_sc_hd__inv_1
XU$$3572 _553_/Q U$$3612/A2 _554_/Q U$$3612/B2 VGND VGND VPWR VPWR U$$3573/A sky130_fd_sc_hd__a22o_1
XFILLER_129_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3583 U$$3583/A U$$3609/B VGND VGND VPWR VPWR U$$3583/X sky130_fd_sc_hd__xor2_1
XFILLER_207_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3594 U$$4140/B1 U$$3636/A2 U$$4007/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3595/A
+ sky130_fd_sc_hd__a22o_1
XU$$2860 _608_/Q U$$2866/A2 _609_/Q U$$2866/B2 VGND VGND VPWR VPWR U$$2861/A sky130_fd_sc_hd__a22o_1
XU$$2871 U$$2871/A _657_/Q VGND VGND VPWR VPWR U$$2871/X sky130_fd_sc_hd__xor2_1
XFILLER_40_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2882 U$$2880/B U$$2877/A _658_/Q U$$2877/Y VGND VGND VPWR VPWR U$$2882/X sky130_fd_sc_hd__a22o_4
XU$$2893 U$$3713/B1 U$$2943/A2 U$$2893/B1 U$$2943/B2 VGND VGND VPWR VPWR U$$2894/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_69_2 dadda_fa_4_69_2/A dadda_fa_4_69_2/B dadda_fa_4_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/CIN dadda_fa_5_69_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_1_36_1 U$$478/X U$$611/X VGND VGND VPWR VPWR dadda_fa_2_37_5/B dadda_fa_3_36_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_102_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_39_0 dadda_fa_7_39_0/A dadda_fa_7_39_0/B dadda_fa_7_39_0/CIN VGND VGND
+ VPWR VPWR _464_/D _335_/D sky130_fd_sc_hd__fa_1
XFILLER_29_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_399 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$705 U$$705/A1 U$$725/A2 U$$707/A1 U$$725/B2 VGND VGND VPWR VPWR U$$706/A sky130_fd_sc_hd__a22o_1
XFILLER_60_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$716 U$$716/A U$$766/B VGND VGND VPWR VPWR U$$716/X sky130_fd_sc_hd__xor2_1
XFILLER_29_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_42_0 U$$91/X U$$224/X U$$357/X VGND VGND VPWR VPWR dadda_fa_2_43_3/A dadda_fa_2_42_4/CIN
+ sky130_fd_sc_hd__fa_1
XU$$727 U$$42/A1 U$$795/A2 U$$42/B1 U$$795/B2 VGND VGND VPWR VPWR U$$728/A sky130_fd_sc_hd__a22o_1
XU$$738 U$$738/A U$$748/B VGND VGND VPWR VPWR U$$738/X sky130_fd_sc_hd__xor2_1
XFILLER_186_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_328 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$749 U$$749/A1 U$$765/A2 U$$749/B1 U$$765/B2 VGND VGND VPWR VPWR U$$750/A sky130_fd_sc_hd__a22o_1
XFILLER_147_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_670 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_336 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1605 U$$3320/A1 VGND VGND VPWR VPWR U$$32/A1 sky130_fd_sc_hd__buf_4
Xrepeater1616 U$$4140/A1 VGND VGND VPWR VPWR U$$3453/B1 sky130_fd_sc_hd__buf_6
XFILLER_137_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1627 _562_/Q VGND VGND VPWR VPWR U$$4273/B1 sky130_fd_sc_hd__buf_6
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1638 U$$3447/B1 VGND VGND VPWR VPWR U$$981/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_153_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1649 U$$2625/A1 VGND VGND VPWR VPWR U$$568/B1 sky130_fd_sc_hd__buf_4
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_76 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_71_2 dadda_fa_3_71_2/A dadda_fa_3_71_2/B dadda_fa_3_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_1/A dadda_fa_4_71_2/B sky130_fd_sc_hd__fa_1
XFILLER_105_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_64_1 dadda_fa_3_64_1/A dadda_fa_3_64_1/B dadda_fa_3_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_0/CIN dadda_fa_4_64_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_41_0 dadda_fa_6_41_0/A dadda_fa_6_41_0/B dadda_fa_6_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_42_0/B dadda_fa_7_41_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_57_0 dadda_fa_3_57_0/A dadda_fa_3_57_0/B dadda_fa_3_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_0/B dadda_fa_4_57_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_43_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2101 U$$2375/A1 U$$2109/A2 U$$2375/B1 U$$2109/B2 VGND VGND VPWR VPWR U$$2102/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2112 U$$2112/A U$$2191/A VGND VGND VPWR VPWR U$$2112/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_100_2 dadda_fa_4_100_2/A dadda_fa_4_100_2/B dadda_fa_4_100_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/CIN dadda_fa_5_100_1/CIN sky130_fd_sc_hd__fa_1
XU$$2123 U$$66/B1 U$$2135/A2 U$$890/B1 U$$2135/B2 VGND VGND VPWR VPWR U$$2124/A sky130_fd_sc_hd__a22o_1
XU$$2134 U$$2134/A U$$2136/B VGND VGND VPWR VPWR U$$2134/X sky130_fd_sc_hd__xor2_1
XU$$1400 U$$715/A1 U$$1428/A2 U$$715/B1 U$$1428/B2 VGND VGND VPWR VPWR U$$1401/A sky130_fd_sc_hd__a22o_1
XU$$2145 U$$2830/A1 U$$2145/A2 U$$229/A1 U$$2145/B2 VGND VGND VPWR VPWR U$$2146/A
+ sky130_fd_sc_hd__a22o_1
XU$$2156 U$$2156/A U$$2191/A VGND VGND VPWR VPWR U$$2156/X sky130_fd_sc_hd__xor2_1
XU$$1411 U$$1411/A U$$1429/B VGND VGND VPWR VPWR U$$1411/X sky130_fd_sc_hd__xor2_1
XU$$1422 U$$463/A1 U$$1458/A2 U$$463/B1 U$$1458/B2 VGND VGND VPWR VPWR U$$1423/A sky130_fd_sc_hd__a22o_1
XU$$2167 U$$2715/A1 U$$2169/A2 U$$525/A1 U$$2169/B2 VGND VGND VPWR VPWR U$$2168/A
+ sky130_fd_sc_hd__a22o_1
XU$$1433 U$$1433/A U$$1479/B VGND VGND VPWR VPWR U$$1433/X sky130_fd_sc_hd__xor2_1
XFILLER_22_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2178 U$$2178/A U$$2186/B VGND VGND VPWR VPWR U$$2178/X sky130_fd_sc_hd__xor2_1
XU$$2189 U$$956/A1 U$$2189/A2 U$$2189/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2190/A
+ sky130_fd_sc_hd__a22o_1
XU$$1444 U$$3088/A1 U$$1486/A2 U$$76/A1 U$$1486/B2 VGND VGND VPWR VPWR U$$1445/A sky130_fd_sc_hd__a22o_1
XFILLER_16_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1455 U$$1455/A U$$1479/B VGND VGND VPWR VPWR U$$1455/X sky130_fd_sc_hd__xor2_1
XFILLER_163_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1466 U$$2971/B1 U$$1474/A2 U$$2838/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1467/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1477 U$$1477/A U$$1507/A VGND VGND VPWR VPWR U$$1477/X sky130_fd_sc_hd__xor2_1
XFILLER_188_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1488 U$$2858/A1 U$$1500/A2 U$$2721/B1 U$$1500/B2 VGND VGND VPWR VPWR U$$1489/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1499 U$$1499/A U$$1501/B VGND VGND VPWR VPWR U$$1499/X sky130_fd_sc_hd__xor2_1
XFILLER_148_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2463_1734 VGND VGND VPWR VPWR U$$2463_1734/HI U$$2463/B1 sky130_fd_sc_hd__conb_1
XFILLER_198_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_114_0 dadda_fa_7_114_0/A dadda_fa_7_114_0/B dadda_fa_7_114_0/CIN VGND
+ VGND VPWR VPWR _539_/D _410_/D sky130_fd_sc_hd__fa_1
XFILLER_50_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_79_1 dadda_fa_5_79_1/A dadda_fa_5_79_1/B dadda_fa_5_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_80_0/B dadda_fa_7_79_0/A sky130_fd_sc_hd__fa_1
XFILLER_83_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$107 _531_/Q _403_/Q VGND VGND VPWR VPWR final_adder.U$$235/B1 final_adder.U$$729/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$118 _542_/Q _414_/Q VGND VGND VPWR VPWR final_adder.U$$613/B1 final_adder.U$$740/A
+ sky130_fd_sc_hd__ha_2
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$129 final_adder.U$$623/A final_adder.U$$623/B final_adder.U$$129/B1
+ VGND VGND VPWR VPWR final_adder.U$$624/B sky130_fd_sc_hd__a21o_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater388 U$$997/A2 VGND VGND VPWR VPWR U$$999/A2 sky130_fd_sc_hd__buf_4
XU$$4070 U$$4070/A U$$4070/B VGND VGND VPWR VPWR U$$4070/X sky130_fd_sc_hd__xor2_1
XFILLER_122_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4081 U$$4490/B1 U$$4095/A2 U$$4357/A1 U$$4081/B2 VGND VGND VPWR VPWR U$$4082/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater399 U$$948/A2 VGND VGND VPWR VPWR U$$956/A2 sky130_fd_sc_hd__buf_6
XU$$4092 U$$4092/A U$$4096/B VGND VGND VPWR VPWR U$$4092/X sky130_fd_sc_hd__xor2_1
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3380 U$$3380/A1 U$$3404/A2 U$$4065/B1 U$$3404/B2 VGND VGND VPWR VPWR U$$3381/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3391 U$$3391/A U$$3397/B VGND VGND VPWR VPWR U$$3391/X sky130_fd_sc_hd__xor2_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2690 U$$2690/A U$$2730/B VGND VGND VPWR VPWR U$$2690/X sky130_fd_sc_hd__xor2_1
XFILLER_34_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_955 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1069 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_870 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_81_1 dadda_fa_4_81_1/A dadda_fa_4_81_1/B dadda_fa_4_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/B dadda_fa_5_81_1/B sky130_fd_sc_hd__fa_1
XFILLER_162_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_74_0 dadda_fa_4_74_0/A dadda_fa_4_74_0/B dadda_fa_4_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/A dadda_fa_5_74_1/A sky130_fd_sc_hd__fa_1
XFILLER_116_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput103 b[44] VGND VGND VPWR VPWR _596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput114 b[54] VGND VGND VPWR VPWR _606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput125 b[6] VGND VGND VPWR VPWR _558_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput136 c[106] VGND VGND VPWR VPWR input136/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput147 c[116] VGND VGND VPWR VPWR input147/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput158 c[126] VGND VGND VPWR VPWR input158/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput169 c[20] VGND VGND VPWR VPWR input169/X sky130_fd_sc_hd__clkbuf_4
Xfinal_adder.U$$630 final_adder.U$$8/SUM final_adder.U$$630/B VGND VGND VPWR VPWR
+ _176_/D sky130_fd_sc_hd__xor2_1
XTAP_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_641_ _642_/CLK _641_/D VGND VGND VPWR VPWR _641_/Q sky130_fd_sc_hd__dfxtp_2
Xfinal_adder.U$$641 final_adder.U$$641/A final_adder.U$$641/B VGND VGND VPWR VPWR
+ _187_/D sky130_fd_sc_hd__xor2_4
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$652 final_adder.U$$652/A final_adder.U$$652/B VGND VGND VPWR VPWR
+ _198_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$663 final_adder.U$$663/A final_adder.U$$663/B VGND VGND VPWR VPWR
+ _209_/D sky130_fd_sc_hd__xor2_2
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$502 U$$502/A U$$518/B VGND VGND VPWR VPWR U$$502/X sky130_fd_sc_hd__xor2_1
XTAP_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$674 final_adder.U$$674/A final_adder.U$$674/B VGND VGND VPWR VPWR
+ _220_/D sky130_fd_sc_hd__xor2_1
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$513 U$$648/B1 U$$517/A2 U$$650/B1 U$$517/B2 VGND VGND VPWR VPWR U$$514/A sky130_fd_sc_hd__a22o_1
XFILLER_45_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$685 final_adder.U$$685/A final_adder.U$$685/B VGND VGND VPWR VPWR
+ _231_/D sky130_fd_sc_hd__xor2_1
XFILLER_186_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$524 U$$524/A U$$547/A VGND VGND VPWR VPWR U$$524/X sky130_fd_sc_hd__xor2_1
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$696 final_adder.U$$696/A final_adder.U$$696/B VGND VGND VPWR VPWR
+ _242_/D sky130_fd_sc_hd__xor2_2
X_572_ _572_/CLK _572_/D VGND VGND VPWR VPWR _572_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$535 U$$944/B1 U$$415/X U$$674/A1 U$$416/X VGND VGND VPWR VPWR U$$536/A sky130_fd_sc_hd__a22o_1
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$546 U$$546/A U$$547/A VGND VGND VPWR VPWR U$$546/X sky130_fd_sc_hd__xor2_1
XFILLER_204_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$557 U$$557/A U$$627/B VGND VGND VPWR VPWR U$$557/X sky130_fd_sc_hd__xor2_1
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$568 U$$705/A1 U$$622/A2 U$$568/B1 U$$622/B2 VGND VGND VPWR VPWR U$$569/A sky130_fd_sc_hd__a22o_1
XU$$579 U$$579/A U$$613/B VGND VGND VPWR VPWR U$$579/X sky130_fd_sc_hd__xor2_1
XFILLER_186_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_89_0 dadda_fa_6_89_0/A dadda_fa_6_89_0/B dadda_fa_6_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_90_0/B dadda_fa_7_89_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1402 _590_/Q VGND VGND VPWR VPWR U$$4468/A1 sky130_fd_sc_hd__buf_4
XFILLER_158_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1413 U$$628/A1 VGND VGND VPWR VPWR U$$491/A1 sky130_fd_sc_hd__buf_8
XFILLER_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1424 U$$3503/A1 VGND VGND VPWR VPWR U$$624/B1 sky130_fd_sc_hd__buf_4
Xrepeater1435 U$$3088/A1 VGND VGND VPWR VPWR U$$74/A1 sky130_fd_sc_hd__buf_4
XFILLER_4_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1446 U$$4317/B1 VGND VGND VPWR VPWR U$$3221/B1 sky130_fd_sc_hd__buf_8
XFILLER_126_778 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1457 U$$4180/A1 VGND VGND VPWR VPWR U$$3769/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1468 U$$749/B1 VGND VGND VPWR VPWR U$$614/A1 sky130_fd_sc_hd__buf_6
XFILLER_207_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1479 U$$4448/A1 VGND VGND VPWR VPWR U$$749/A1 sky130_fd_sc_hd__buf_6
XFILLER_119_1139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1230 U$$817/B1 U$$1230/A2 U$$1230/B1 U$$1230/B2 VGND VGND VPWR VPWR U$$1231/A
+ sky130_fd_sc_hd__a22o_1
XU$$1241 U$$828/B1 U$$1295/A2 U$$556/B1 U$$1295/B2 VGND VGND VPWR VPWR U$$1242/A sky130_fd_sc_hd__a22o_1
XU$$1252 U$$1252/A U$$1296/B VGND VGND VPWR VPWR U$$1252/X sky130_fd_sc_hd__xor2_1
XFILLER_188_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1263 U$$989/A1 U$$1291/A2 U$$32/A1 U$$1291/B2 VGND VGND VPWR VPWR U$$1264/A sky130_fd_sc_hd__a22o_1
XU$$1274 U$$1274/A U$$1280/B VGND VGND VPWR VPWR U$$1274/X sky130_fd_sc_hd__xor2_1
XFILLER_188_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1285 U$$463/A1 U$$1291/A2 U$$463/B1 U$$1291/B2 VGND VGND VPWR VPWR U$$1286/A sky130_fd_sc_hd__a22o_1
XFILLER_203_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1296 U$$1296/A U$$1296/B VGND VGND VPWR VPWR U$$1296/X sky130_fd_sc_hd__xor2_1
XFILLER_188_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_91_0 dadda_fa_5_91_0/A dadda_fa_5_91_0/B dadda_fa_5_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_92_0/A dadda_fa_6_91_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_190_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_76_6 U$$3883/X U$$4016/X U$$4149/X VGND VGND VPWR VPWR dadda_fa_2_77_2/B
+ dadda_fa_2_76_5/B sky130_fd_sc_hd__fa_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_5 U$$4401/X input222/X dadda_fa_1_69_5/CIN VGND VGND VPWR VPWR dadda_fa_2_70_2/A
+ dadda_fa_2_69_5/A sky130_fd_sc_hd__fa_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_96_0 dadda_ha_1_96_0/A U$$2327/X VGND VGND VPWR VPWR dadda_fa_3_97_0/A
+ dadda_fa_3_96_0/A sky130_fd_sc_hd__ha_1
XFILLER_10_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_100_1 dadda_fa_3_100_1/A dadda_fa_3_100_1/B dadda_fa_3_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_0/CIN dadda_fa_4_100_2/A sky130_fd_sc_hd__fa_1
XFILLER_101_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_121_0 dadda_fa_6_121_0/A dadda_fa_6_121_0/B dadda_fa_6_121_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_122_0/B dadda_fa_7_121_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_64_4 U$$1731/X U$$1864/X U$$1997/X VGND VGND VPWR VPWR dadda_fa_1_65_6/CIN
+ dadda_fa_1_64_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_41_3 dadda_fa_3_41_3/A dadda_fa_3_41_3/B dadda_fa_3_41_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_1/B dadda_fa_4_41_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_97_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$471 final_adder.U$$294/B final_adder.U$$698/B final_adder.U$$205/X
+ VGND VGND VPWR VPWR final_adder.U$$700/B sky130_fd_sc_hd__a21o_1
XTAP_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$310 U$$310/A1 U$$318/A2 U$$449/A1 U$$318/B2 VGND VGND VPWR VPWR U$$311/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_34_2 dadda_fa_3_34_2/A dadda_fa_3_34_2/B dadda_fa_3_34_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_1/A dadda_fa_4_34_2/B sky130_fd_sc_hd__fa_1
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_624_ _624_/CLK _624_/D VGND VGND VPWR VPWR _624_/Q sky130_fd_sc_hd__dfxtp_1
XU$$321 U$$321/A U$$335/B VGND VGND VPWR VPWR U$$321/X sky130_fd_sc_hd__xor2_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$332 U$$58/A1 U$$398/A2 U$$60/A1 U$$398/B2 VGND VGND VPWR VPWR U$$333/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$493 final_adder.U$$316/B final_adder.U$$742/B final_adder.U$$249/X
+ VGND VGND VPWR VPWR final_adder.U$$744/B sky130_fd_sc_hd__a21o_1
XFILLER_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$343 U$$343/A U$$351/B VGND VGND VPWR VPWR U$$343/X sky130_fd_sc_hd__xor2_1
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$354 U$$491/A1 U$$398/A2 U$$493/A1 U$$398/B2 VGND VGND VPWR VPWR U$$355/A sky130_fd_sc_hd__a22o_1
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_27_1 U$$1524/X U$$1657/X U$$1790/X VGND VGND VPWR VPWR dadda_fa_4_28_0/CIN
+ dadda_fa_4_27_2/A sky130_fd_sc_hd__fa_1
XFILLER_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$365 U$$365/A U$$410/A VGND VGND VPWR VPWR U$$365/X sky130_fd_sc_hd__xor2_1
X_555_ _558_/CLK _555_/D VGND VGND VPWR VPWR _555_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$376 U$$648/B1 U$$384/A2 U$$650/B1 U$$384/B2 VGND VGND VPWR VPWR U$$377/A sky130_fd_sc_hd__a22o_1
XFILLER_60_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$387 U$$387/A U$$393/B VGND VGND VPWR VPWR U$$387/X sky130_fd_sc_hd__xor2_1
XU$$398 U$$944/B1 U$$398/A2 U$$674/A1 U$$398/B2 VGND VGND VPWR VPWR U$$399/A sky130_fd_sc_hd__a22o_1
XFILLER_72_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_486_ _486_/CLK _486_/D VGND VGND VPWR VPWR _486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1210 U$$3418/A1 VGND VGND VPWR VPWR U$$4238/B1 sky130_fd_sc_hd__buf_4
Xrepeater1221 U$$3005/A1 VGND VGND VPWR VPWR U$$3551/B1 sky130_fd_sc_hd__buf_4
Xrepeater1232 _610_/Q VGND VGND VPWR VPWR U$$2588/B1 sky130_fd_sc_hd__buf_6
XFILLER_160_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1243 U$$4369/A1 VGND VGND VPWR VPWR U$$805/B1 sky130_fd_sc_hd__buf_4
Xrepeater1254 U$$3269/B1 VGND VGND VPWR VPWR U$$3132/B1 sky130_fd_sc_hd__buf_6
XFILLER_99_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1265 U$$2991/B1 VGND VGND VPWR VPWR U$$251/B1 sky130_fd_sc_hd__buf_6
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_86_5 dadda_fa_2_86_5/A dadda_fa_2_86_5/B dadda_fa_2_86_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_2/A dadda_fa_4_86_0/A sky130_fd_sc_hd__fa_2
Xrepeater1276 U$$4498/A1 VGND VGND VPWR VPWR U$$936/A1 sky130_fd_sc_hd__buf_4
XFILLER_114_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1287 U$$3674/A1 VGND VGND VPWR VPWR U$$4222/A1 sky130_fd_sc_hd__buf_4
XFILLER_113_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1298 U$$3122/A1 VGND VGND VPWR VPWR U$$517/B1 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_2_79_4 dadda_fa_2_79_4/A dadda_fa_2_79_4/B dadda_fa_2_79_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/CIN dadda_fa_3_79_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_171_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1060 U$$1060/A U$$996/B VGND VGND VPWR VPWR U$$1060/X sky130_fd_sc_hd__xor2_1
XFILLER_189_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1071 U$$934/A1 U$$963/X U$$936/A1 U$$964/X VGND VGND VPWR VPWR U$$1072/A sky130_fd_sc_hd__a22o_1
XFILLER_51_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1082 U$$1082/A U$$1095/A VGND VGND VPWR VPWR U$$1082/X sky130_fd_sc_hd__xor2_1
XFILLER_32_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1093 U$$956/A1 U$$1093/A2 U$$1093/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1094/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_116_1 dadda_fa_5_116_1/A dadda_fa_5_116_1/B dadda_fa_5_116_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_117_0/B dadda_fa_7_116_0/A sky130_fd_sc_hd__fa_1
XFILLER_136_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_109_0 dadda_fa_5_109_0/A dadda_fa_5_109_0/B dadda_fa_5_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_110_0/A dadda_fa_6_109_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_81_4 U$$2829/X U$$2962/X U$$3095/X VGND VGND VPWR VPWR dadda_fa_2_82_2/B
+ dadda_fa_2_81_5/A sky130_fd_sc_hd__fa_1
XFILLER_208_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_74_3 U$$2948/X U$$3081/X U$$3214/X VGND VGND VPWR VPWR dadda_fa_2_75_1/B
+ dadda_fa_2_74_4/B sky130_fd_sc_hd__fa_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_51_2 dadda_fa_4_51_2/A dadda_fa_4_51_2/B dadda_fa_4_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/CIN dadda_fa_5_51_1/CIN sky130_fd_sc_hd__fa_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_2 U$$3333/X U$$3466/X U$$3599/X VGND VGND VPWR VPWR dadda_fa_2_68_1/A
+ dadda_fa_2_67_4/A sky130_fd_sc_hd__fa_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_44_1 dadda_fa_4_44_1/A dadda_fa_4_44_1/B dadda_fa_4_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/B dadda_fa_5_44_1/B sky130_fd_sc_hd__fa_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_21_0 dadda_fa_7_21_0/A dadda_fa_7_21_0/B dadda_fa_7_21_0/CIN VGND VGND
+ VPWR VPWR _446_/D _317_/D sky130_fd_sc_hd__fa_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_37_0 dadda_fa_4_37_0/A dadda_fa_4_37_0/B dadda_fa_4_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/A dadda_fa_5_37_1/A sky130_fd_sc_hd__fa_1
XFILLER_73_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ _455_/CLK _340_/D VGND VGND VPWR VPWR _340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_271_ _521_/CLK _271_/D VGND VGND VPWR VPWR _271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_0_70_4 U$$2009/X U$$2142/X VGND VGND VPWR VPWR dadda_fa_1_71_7/CIN dadda_fa_2_70_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_68_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_89_3 dadda_fa_3_89_3/A dadda_fa_3_89_3/B dadda_fa_3_89_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_1/B dadda_fa_4_89_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_56_2 U$$917/X U$$1050/X VGND VGND VPWR VPWR dadda_fa_1_57_8/A dadda_fa_2_56_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_2_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_62_1 U$$530/X U$$663/X U$$796/X VGND VGND VPWR VPWR dadda_fa_1_63_5/CIN
+ dadda_fa_1_62_7/CIN sky130_fd_sc_hd__fa_1
XU$$3696_1754 VGND VGND VPWR VPWR U$$3696_1754/HI U$$3696/B1 sky130_fd_sc_hd__conb_1
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3902 U$$3902/A1 U$$3958/A2 U$$3902/B1 U$$3958/B2 VGND VGND VPWR VPWR U$$3903/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_55_0 U$$117/X U$$250/X U$$383/X VGND VGND VPWR VPWR dadda_fa_1_56_7/CIN
+ dadda_fa_1_55_8/CIN sky130_fd_sc_hd__fa_1
XU$$3913 U$$3913/A U$$3933/B VGND VGND VPWR VPWR U$$3913/X sky130_fd_sc_hd__xor2_1
XFILLER_91_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3924 _592_/Q U$$3932/A2 _593_/Q U$$3932/B2 VGND VGND VPWR VPWR U$$3925/A sky130_fd_sc_hd__a22o_1
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3935 U$$3935/A U$$3935/B VGND VGND VPWR VPWR U$$3935/X sky130_fd_sc_hd__xor2_1
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3946 U$$4355/B1 U$$3968/A2 U$$4222/A1 U$$3968/B2 VGND VGND VPWR VPWR U$$3947/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3957 U$$3957/A U$$3965/B VGND VGND VPWR VPWR U$$3957/X sky130_fd_sc_hd__xor2_1
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$290 final_adder.U$$290/A final_adder.U$$290/B VGND VGND VPWR VPWR
+ final_adder.U$$336/A sky130_fd_sc_hd__and2_1
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3968 U$$4516/A1 U$$3968/A2 U$$4516/B1 U$$3968/B2 VGND VGND VPWR VPWR U$$3969/A
+ sky130_fd_sc_hd__a22o_1
XU$$140 U$$272/B U$$140/B VGND VGND VPWR VPWR U$$140/X sky130_fd_sc_hd__and2_1
XFILLER_91_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_607_ _613_/CLK _607_/D VGND VGND VPWR VPWR _607_/Q sky130_fd_sc_hd__dfxtp_1
XU$$151 U$$14/A1 U$$181/A2 U$$16/A1 U$$181/B2 VGND VGND VPWR VPWR U$$152/A sky130_fd_sc_hd__a22o_1
XFILLER_79_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3979 U$$3979/A1 U$$4005/A2 U$$4392/A1 U$$4005/B2 VGND VGND VPWR VPWR U$$3980/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$162 U$$162/A U$$190/B VGND VGND VPWR VPWR U$$162/X sky130_fd_sc_hd__xor2_1
XFILLER_150_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$173 U$$36/A1 U$$195/A2 U$$38/A1 U$$195/B2 VGND VGND VPWR VPWR U$$174/A sky130_fd_sc_hd__a22o_1
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$184 U$$184/A U$$232/B VGND VGND VPWR VPWR U$$184/X sky130_fd_sc_hd__xor2_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$195 U$$58/A1 U$$195/A2 U$$60/A1 U$$195/B2 VGND VGND VPWR VPWR U$$196/A sky130_fd_sc_hd__a22o_1
XFILLER_72_392 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_538_ _538_/CLK _538_/D VGND VGND VPWR VPWR _538_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_469_ _469_/CLK _469_/D VGND VGND VPWR VPWR _469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_91_3 U$$4312/X U$$4445/X input247/X VGND VGND VPWR VPWR dadda_fa_3_92_1/B
+ dadda_fa_3_91_3/B sky130_fd_sc_hd__fa_1
XFILLER_142_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1040 U$$2303/B VGND VGND VPWR VPWR U$$2243/B sky130_fd_sc_hd__buf_6
XFILLER_173_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1051 U$$2170/B VGND VGND VPWR VPWR U$$2144/B sky130_fd_sc_hd__buf_8
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1062 U$$2043/B VGND VGND VPWR VPWR U$$2054/A sky130_fd_sc_hd__buf_6
Xdadda_fa_2_84_2 dadda_fa_2_84_2/A dadda_fa_2_84_2/B dadda_fa_2_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/A dadda_fa_3_84_3/A sky130_fd_sc_hd__fa_1
Xoutput259 _269_/Q VGND VGND VPWR VPWR o[101] sky130_fd_sc_hd__buf_2
Xrepeater1073 _643_/Q VGND VGND VPWR VPWR U$$1918/A sky130_fd_sc_hd__buf_4
Xrepeater1084 U$$1598/B VGND VGND VPWR VPWR U$$1554/B sky130_fd_sc_hd__buf_6
Xrepeater1095 U$$1479/B VGND VGND VPWR VPWR U$$1443/B sky130_fd_sc_hd__buf_6
Xdadda_fa_5_61_1 dadda_fa_5_61_1/A dadda_fa_5_61_1/B dadda_fa_5_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_62_0/B dadda_fa_7_61_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_77_1 dadda_fa_2_77_1/A dadda_fa_2_77_1/B dadda_fa_2_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_0/CIN dadda_fa_3_77_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_173_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_54_0 dadda_fa_5_54_0/A dadda_fa_5_54_0/B dadda_fa_5_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_55_0/A dadda_fa_6_54_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_8 U$$3571/X input205/X dadda_fa_1_53_8/CIN VGND VGND VPWR VPWR dadda_fa_2_54_3/A
+ dadda_fa_3_53_0/A sky130_fd_sc_hd__fa_1
XFILLER_68_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_100_0 dadda_fa_2_100_0/A U$$2601/X U$$2734/X VGND VGND VPWR VPWR dadda_fa_3_101_1/B
+ dadda_fa_3_100_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_51_532 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_99_2 dadda_fa_4_99_2/A dadda_fa_4_99_2/B dadda_fa_4_99_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/CIN dadda_fa_5_99_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_165_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_692 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_69_0 dadda_fa_7_69_0/A dadda_fa_7_69_0/B dadda_fa_7_69_0/CIN VGND VGND
+ VPWR VPWR _494_/D _365_/D sky130_fd_sc_hd__fa_1
XFILLER_117_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_72_0 U$$2013/X U$$2146/X U$$2279/X VGND VGND VPWR VPWR dadda_fa_2_73_0/B
+ dadda_fa_2_72_3/B sky130_fd_sc_hd__fa_1
XFILLER_59_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1014 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3209 U$$467/B1 U$$3209/A2 U$$4031/B1 U$$3209/B2 VGND VGND VPWR VPWR U$$3210/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2508 U$$2508/A1 U$$2550/A2 U$$2508/B1 U$$2550/B2 VGND VGND VPWR VPWR U$$2509/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2519 U$$2519/A U$$2541/B VGND VGND VPWR VPWR U$$2519/X sky130_fd_sc_hd__xor2_1
XFILLER_15_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1807 U$$4410/A1 U$$1843/A2 U$$3042/A1 U$$1843/B2 VGND VGND VPWR VPWR U$$1808/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1818 U$$1818/A U$$1820/B VGND VGND VPWR VPWR U$$1818/X sky130_fd_sc_hd__xor2_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1829 U$$4158/A1 U$$1855/A2 U$$50/A1 U$$1855/B2 VGND VGND VPWR VPWR U$$1830/A sky130_fd_sc_hd__a22o_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_323_ _451_/CLK _323_/D VGND VGND VPWR VPWR _323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_254_ _379_/CLK _254_/D VGND VGND VPWR VPWR _254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_784 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_934 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_185_ _189_/CLK _185_/D VGND VGND VPWR VPWR _185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_94_1 dadda_fa_3_94_1/A dadda_fa_3_94_1/B dadda_fa_3_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_0/CIN dadda_fa_4_94_2/A sky130_fd_sc_hd__fa_1
XFILLER_155_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_71_0 dadda_fa_6_71_0/A dadda_fa_6_71_0/B dadda_fa_6_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_72_0/B dadda_fa_7_71_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_87_0 dadda_fa_3_87_0/A dadda_fa_3_87_0/B dadda_fa_3_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_0/B dadda_fa_4_87_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater707 U$$3958/B2 VGND VGND VPWR VPWR U$$3970/B2 sky130_fd_sc_hd__buf_4
XU$$4400 U$$4400/A1 U$$4388/X U$$4402/A1 U$$4438/B2 VGND VGND VPWR VPWR U$$4401/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater718 U$$3628/B2 VGND VGND VPWR VPWR U$$3612/B2 sky130_fd_sc_hd__buf_6
XU$$4411 U$$4411/A U$$4411/B VGND VGND VPWR VPWR U$$4411/X sky130_fd_sc_hd__xor2_1
Xrepeater729 U$$3537/B2 VGND VGND VPWR VPWR U$$3531/B2 sky130_fd_sc_hd__buf_4
XFILLER_133_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4422 _567_/Q U$$4388/X _568_/Q U$$4454/B2 VGND VGND VPWR VPWR U$$4423/A sky130_fd_sc_hd__a22o_1
XU$$4433 U$$4433/A U$$4433/B VGND VGND VPWR VPWR U$$4433/X sky130_fd_sc_hd__xor2_1
XU$$4444 U$$4444/A1 U$$4388/X U$$4444/B1 U$$4480/B2 VGND VGND VPWR VPWR U$$4445/A
+ sky130_fd_sc_hd__a22o_1
XU$$4455 U$$4455/A U$$4455/B VGND VGND VPWR VPWR U$$4455/X sky130_fd_sc_hd__xor2_2
XU$$3710 U$$3710/A U$$3764/B VGND VGND VPWR VPWR U$$3710/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_49_5 dadda_fa_2_49_5/A dadda_fa_2_49_5/B dadda_fa_2_49_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_2/A dadda_fa_4_49_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_116_0 U$$3830/X U$$3963/X U$$4096/X VGND VGND VPWR VPWR dadda_fa_5_117_0/A
+ dadda_fa_5_116_1/A sky130_fd_sc_hd__fa_1
XFILLER_37_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3721 U$$4269/A1 U$$3769/A2 U$$4408/A1 U$$3769/B2 VGND VGND VPWR VPWR U$$3722/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4466 U$$4466/A1 U$$4388/X U$$4468/A1 U$$4468/B2 VGND VGND VPWR VPWR U$$4467/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3732 U$$3732/A U$$3816/B VGND VGND VPWR VPWR U$$3732/X sky130_fd_sc_hd__xor2_1
XU$$4477 U$$4477/A U$$4477/B VGND VGND VPWR VPWR U$$4477/X sky130_fd_sc_hd__xor2_1
XFILLER_93_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4488 U$$926/A1 U$$4388/X U$$928/A1 U$$4496/B2 VGND VGND VPWR VPWR U$$4489/A sky130_fd_sc_hd__a22o_1
XFILLER_18_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3743 U$$4291/A1 U$$3743/A2 U$$4293/A1 U$$3743/B2 VGND VGND VPWR VPWR U$$3744/A
+ sky130_fd_sc_hd__a22o_1
XU$$3754 U$$3754/A U$$3800/B VGND VGND VPWR VPWR U$$3754/X sky130_fd_sc_hd__xor2_1
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4499 U$$4499/A U$$4499/B VGND VGND VPWR VPWR U$$4499/X sky130_fd_sc_hd__xor2_1
XFILLER_18_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3765 U$$4176/A1 U$$3777/A2 U$$4176/B1 U$$3777/B2 VGND VGND VPWR VPWR U$$3766/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3776 U$$3776/A _671_/Q VGND VGND VPWR VPWR U$$3776/X sky130_fd_sc_hd__xor2_1
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3787 U$$4061/A1 U$$3795/A2 _593_/Q U$$3795/B2 VGND VGND VPWR VPWR U$$3788/A sky130_fd_sc_hd__a22o_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3798 U$$3798/A U$$3804/B VGND VGND VPWR VPWR U$$3798/X sky130_fd_sc_hd__xor2_1
XFILLER_79_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_380 U$$922/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_391 U$$1478/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_51_5 U$$2104/X U$$2237/X U$$2370/X VGND VGND VPWR VPWR dadda_fa_2_52_2/A
+ dadda_fa_2_51_5/A sky130_fd_sc_hd__fa_1
XU$$909 U$$909/A U$$958/A VGND VGND VPWR VPWR U$$909/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_44_4 U$$1691/X U$$1824/X U$$1957/X VGND VGND VPWR VPWR dadda_fa_2_45_3/CIN
+ dadda_fa_2_44_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_14_2 U$$994/B input162/X dadda_ha_3_14_0/SUM VGND VGND VPWR VPWR dadda_fa_5_15_0/CIN
+ dadda_fa_5_14_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_34_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_78_0_1873 VGND VGND VPWR VPWR dadda_ha_0_78_0/A dadda_ha_0_78_0_1873/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_24_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_727 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4489_1823 VGND VGND VPWR VPWR U$$4489_1823/HI U$$4489/B sky130_fd_sc_hd__conb_1
XFILLER_59_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3006 U$$3006/A U$$3008/B VGND VGND VPWR VPWR U$$3006/X sky130_fd_sc_hd__xor2_1
XFILLER_207_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3017 _661_/Q U$$3017/B VGND VGND VPWR VPWR U$$3017/X sky130_fd_sc_hd__and2_1
XU$$3028 U$$3163/B1 U$$3054/A2 U$$3713/B1 U$$3054/B2 VGND VGND VPWR VPWR U$$3029/A
+ sky130_fd_sc_hd__a22o_1
XU$$3039 U$$3039/A U$$3049/B VGND VGND VPWR VPWR U$$3039/X sky130_fd_sc_hd__xor2_1
XU$$2305 U$$2305/A U$$2309/B VGND VGND VPWR VPWR U$$2305/X sky130_fd_sc_hd__xor2_1
XU$$2316 U$$2999/B1 U$$2318/A2 U$$946/B1 U$$2318/B2 VGND VGND VPWR VPWR U$$2317/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2327 U$$2327/A U$$2328/A VGND VGND VPWR VPWR U$$2327/X sky130_fd_sc_hd__xor2_1
XU$$2338 U$$2338/A U$$2418/B VGND VGND VPWR VPWR U$$2338/X sky130_fd_sc_hd__xor2_1
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1604 U$$1604/A U$$1642/B VGND VGND VPWR VPWR U$$1604/X sky130_fd_sc_hd__xor2_1
XU$$2349 U$$840/B1 U$$2395/A2 U$$2625/A1 U$$2395/B2 VGND VGND VPWR VPWR U$$2350/A
+ sky130_fd_sc_hd__a22o_1
XU$$1615 U$$2983/B1 U$$1635/A2 U$$2848/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1616/A
+ sky130_fd_sc_hd__a22o_1
XU$$1626 U$$1626/A U$$1628/B VGND VGND VPWR VPWR U$$1626/X sky130_fd_sc_hd__xor2_1
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1637 U$$3418/A1 U$$1511/X U$$678/B1 U$$1512/X VGND VGND VPWR VPWR U$$1638/A sky130_fd_sc_hd__a22o_1
XFILLER_163_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1648 U$$1646/Y _640_/Q _639_/Q U$$1647/X U$$1644/Y VGND VGND VPWR VPWR U$$1648/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_72_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1659 U$$1659/A U$$1687/B VGND VGND VPWR VPWR U$$1659/X sky130_fd_sc_hd__xor2_1
XFILLER_72_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_699 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_306_ _435_/CLK _306_/D VGND VGND VPWR VPWR _306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_237_ _503_/CLK _237_/D VGND VGND VPWR VPWR _237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_168_ _179_/CLK _168_/D VGND VGND VPWR VPWR _168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_61_4 dadda_fa_2_61_4/A dadda_fa_2_61_4/B dadda_fa_2_61_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/CIN dadda_fa_3_61_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater504 U$$3082/A2 VGND VGND VPWR VPWR U$$3046/A2 sky130_fd_sc_hd__buf_6
XFILLER_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater515 U$$3005/A2 VGND VGND VPWR VPWR U$$2997/A2 sky130_fd_sc_hd__buf_4
XFILLER_46_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater526 U$$278/X VGND VGND VPWR VPWR U$$408/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_38_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_54_3 dadda_fa_2_54_3/A dadda_fa_2_54_3/B dadda_fa_2_54_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/B dadda_fa_3_54_3/B sky130_fd_sc_hd__fa_1
Xrepeater537 U$$2705/A2 VGND VGND VPWR VPWR U$$2663/A2 sky130_fd_sc_hd__buf_4
XFILLER_78_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater548 U$$2588/A2 VGND VGND VPWR VPWR U$$2600/A2 sky130_fd_sc_hd__buf_6
XU$$4230 U$$805/A1 U$$4238/A2 U$$805/B1 U$$4238/B2 VGND VGND VPWR VPWR U$$4231/A sky130_fd_sc_hd__a22o_1
Xrepeater559 U$$2274/A2 VGND VGND VPWR VPWR U$$2262/A2 sky130_fd_sc_hd__buf_4
XFILLER_77_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4241 U$$4241/A U$$4246/A VGND VGND VPWR VPWR U$$4241/X sky130_fd_sc_hd__xor2_1
XFILLER_93_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4252 U$$4250/B U$$4203/B _678_/Q U$$4247/Y VGND VGND VPWR VPWR U$$4252/X sky130_fd_sc_hd__a22o_1
XU$$4263 _556_/Q U$$4347/A2 U$$4402/A1 U$$4347/B2 VGND VGND VPWR VPWR U$$4264/A sky130_fd_sc_hd__a22o_1
XFILLER_38_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_47_2 dadda_fa_2_47_2/A dadda_fa_2_47_2/B dadda_fa_2_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/A dadda_fa_3_47_3/A sky130_fd_sc_hd__fa_1
XFILLER_168_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4274 U$$4274/A U$$4296/B VGND VGND VPWR VPWR U$$4274/X sky130_fd_sc_hd__xor2_1
XU$$4285 U$$4285/A1 U$$4327/A2 _568_/Q U$$4319/B2 VGND VGND VPWR VPWR U$$4286/A sky130_fd_sc_hd__a22o_1
XFILLER_66_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3540 U$$3540/A U$$3562/A VGND VGND VPWR VPWR U$$3540/X sky130_fd_sc_hd__xor2_1
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3551 U$$4510/A1 U$$3555/A2 U$$3551/B1 U$$3555/B2 VGND VGND VPWR VPWR U$$3552/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_24_1 dadda_fa_5_24_1/A dadda_fa_5_24_1/B dadda_fa_5_24_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_25_0/B dadda_fa_7_24_0/A sky130_fd_sc_hd__fa_1
XFILLER_207_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4296 U$$4296/A U$$4296/B VGND VGND VPWR VPWR U$$4296/X sky130_fd_sc_hd__xor2_1
XFILLER_53_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3562 U$$3562/A VGND VGND VPWR VPWR U$$3562/Y sky130_fd_sc_hd__inv_1
XU$$3573 U$$3573/A U$$3613/B VGND VGND VPWR VPWR U$$3573/X sky130_fd_sc_hd__xor2_1
XFILLER_209_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_17_0 dadda_fa_5_17_0/A dadda_fa_5_17_0/B dadda_fa_5_17_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_18_0/A dadda_fa_6_17_0/CIN sky130_fd_sc_hd__fa_1
XU$$3584 U$$4404/B1 U$$3628/A2 U$$3584/B1 U$$3628/B2 VGND VGND VPWR VPWR U$$3585/A
+ sky130_fd_sc_hd__a22o_1
XU$$2850 _603_/Q U$$2866/A2 U$$3674/A1 U$$2866/B2 VGND VGND VPWR VPWR U$$2851/A sky130_fd_sc_hd__a22o_1
XU$$3595 U$$3595/A U$$3637/B VGND VGND VPWR VPWR U$$3595/X sky130_fd_sc_hd__xor2_1
XFILLER_197_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2861 U$$2861/A U$$2861/B VGND VGND VPWR VPWR U$$2861/X sky130_fd_sc_hd__xor2_1
XU$$2872 _614_/Q U$$2874/A2 U$$2872/B1 U$$2874/B2 VGND VGND VPWR VPWR U$$2873/A sky130_fd_sc_hd__a22o_1
XU$$2883 U$$2883/A1 U$$2929/A2 U$$3157/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2884/A
+ sky130_fd_sc_hd__a22o_1
XU$$2894 U$$2894/A U$$2944/B VGND VGND VPWR VPWR U$$2894/X sky130_fd_sc_hd__xor2_1
XFILLER_60_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$706 U$$706/A U$$726/B VGND VGND VPWR VPWR U$$706/X sky130_fd_sc_hd__xor2_1
XFILLER_99_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$717 U$$854/A1 U$$759/A2 U$$993/A1 U$$759/B2 VGND VGND VPWR VPWR U$$718/A sky130_fd_sc_hd__a22o_1
XFILLER_186_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_42_1 U$$490/X U$$623/X U$$756/X VGND VGND VPWR VPWR dadda_fa_2_43_3/B
+ dadda_fa_2_42_5/A sky130_fd_sc_hd__fa_1
XU$$728 U$$728/A U$$796/B VGND VGND VPWR VPWR U$$728/X sky130_fd_sc_hd__xor2_1
XFILLER_84_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$739 U$$876/A1 U$$747/A2 U$$878/A1 U$$747/B2 VGND VGND VPWR VPWR U$$740/A sky130_fd_sc_hd__a22o_1
XFILLER_204_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1606 U$$3320/A1 VGND VGND VPWR VPWR U$$854/A1 sky130_fd_sc_hd__buf_6
Xrepeater1617 U$$4140/A1 VGND VGND VPWR VPWR U$$4003/A1 sky130_fd_sc_hd__buf_6
Xrepeater1628 U$$3312/B1 VGND VGND VPWR VPWR U$$848/A1 sky130_fd_sc_hd__buf_6
Xrepeater1639 U$$24/A1 VGND VGND VPWR VPWR U$$22/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_180_543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_71_3 dadda_fa_3_71_3/A dadda_fa_3_71_3/B dadda_fa_3_71_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_1/B dadda_fa_4_71_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_64_2 dadda_fa_3_64_2/A dadda_fa_3_64_2/B dadda_fa_3_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_1/A dadda_fa_4_64_2/B sky130_fd_sc_hd__fa_1
XFILLER_0_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_57_1 dadda_fa_3_57_1/A dadda_fa_3_57_1/B dadda_fa_3_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_0/CIN dadda_fa_4_57_2/A sky130_fd_sc_hd__fa_1
XFILLER_86_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_34_0 dadda_fa_6_34_0/A dadda_fa_6_34_0/B dadda_fa_6_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_35_0/B dadda_fa_7_34_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_120_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2102 U$$2102/A U$$2110/B VGND VGND VPWR VPWR U$$2102/X sky130_fd_sc_hd__xor2_1
XU$$2113 U$$3346/A1 U$$2169/A2 _578_/Q U$$2169/B2 VGND VGND VPWR VPWR U$$2114/A sky130_fd_sc_hd__a22o_1
XFILLER_142_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2124 U$$2124/A U$$2136/B VGND VGND VPWR VPWR U$$2124/X sky130_fd_sc_hd__xor2_1
XU$$2135 U$$3642/A1 U$$2135/A2 U$$3505/B1 U$$2135/B2 VGND VGND VPWR VPWR U$$2136/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1401 U$$1401/A U$$1429/B VGND VGND VPWR VPWR U$$1401/X sky130_fd_sc_hd__xor2_1
XFILLER_62_446 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2146 U$$2146/A U$$2170/B VGND VGND VPWR VPWR U$$2146/X sky130_fd_sc_hd__xor2_1
XU$$2157 U$$3388/B1 U$$2189/A2 U$$3253/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2158/A
+ sky130_fd_sc_hd__a22o_1
XU$$1412 U$$316/A1 U$$1428/A2 U$$44/A1 U$$1428/B2 VGND VGND VPWR VPWR U$$1413/A sky130_fd_sc_hd__a22o_1
XFILLER_90_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1423 U$$1423/A U$$1459/B VGND VGND VPWR VPWR U$$1423/X sky130_fd_sc_hd__xor2_1
XFILLER_50_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2168 U$$2168/A U$$2170/B VGND VGND VPWR VPWR U$$2168/X sky130_fd_sc_hd__xor2_1
XU$$1434 U$$749/A1 U$$1442/A2 U$$614/A1 U$$1442/B2 VGND VGND VPWR VPWR U$$1435/A sky130_fd_sc_hd__a22o_1
XU$$2179 U$$2314/B1 U$$2185/A2 U$$946/B1 U$$2185/B2 VGND VGND VPWR VPWR U$$2180/A
+ sky130_fd_sc_hd__a22o_1
XU$$1445 U$$1445/A U$$1487/B VGND VGND VPWR VPWR U$$1445/X sky130_fd_sc_hd__xor2_1
XFILLER_90_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1456 U$$84/B1 U$$1458/A2 U$$634/B1 U$$1458/B2 VGND VGND VPWR VPWR U$$1457/A sky130_fd_sc_hd__a22o_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1467 U$$1467/A U$$1475/B VGND VGND VPWR VPWR U$$1467/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1478 U$$791/B1 U$$1478/A2 U$$2848/B1 U$$1478/B2 VGND VGND VPWR VPWR U$$1479/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1489 U$$1489/A U$$1501/B VGND VGND VPWR VPWR U$$1489/X sky130_fd_sc_hd__xor2_1
XFILLER_188_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1098 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_107_0 dadda_fa_7_107_0/A dadda_fa_7_107_0/B dadda_fa_7_107_0/CIN VGND
+ VGND VPWR VPWR _532_/D _403_/D sky130_fd_sc_hd__fa_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$108 _532_/Q _404_/Q VGND VGND VPWR VPWR final_adder.U$$603/B1 final_adder.U$$730/A
+ sky130_fd_sc_hd__ha_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$119 _543_/Q _415_/Q VGND VGND VPWR VPWR final_adder.U$$247/B1 final_adder.U$$741/A
+ sky130_fd_sc_hd__ha_2
Xdadda_fa_2_52_0 dadda_fa_2_52_0/A dadda_fa_2_52_0/B dadda_fa_2_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_0/B dadda_fa_3_52_2/B sky130_fd_sc_hd__fa_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3422_1750 VGND VGND VPWR VPWR U$$3422_1750/HI U$$3422/B1 sky130_fd_sc_hd__conb_1
XFILLER_26_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4060 U$$4060/A U$$4070/B VGND VGND VPWR VPWR U$$4060/X sky130_fd_sc_hd__xor2_1
Xrepeater389 U$$963/X VGND VGND VPWR VPWR U$$997/A2 sky130_fd_sc_hd__buf_6
XFILLER_65_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4071 U$$4206/B1 U$$4071/A2 U$$4208/B1 U$$4071/B2 VGND VGND VPWR VPWR U$$4072/A
+ sky130_fd_sc_hd__a22o_1
XU$$4082 U$$4082/A U$$4096/B VGND VGND VPWR VPWR U$$4082/X sky130_fd_sc_hd__xor2_1
XU$$4093 U$$4228/B1 U$$4095/A2 U$$4369/A1 U$$4105/B2 VGND VGND VPWR VPWR U$$4094/A
+ sky130_fd_sc_hd__a22o_1
XU$$3370 U$$3505/B1 U$$3418/A2 U$$3372/A1 U$$3418/B2 VGND VGND VPWR VPWR U$$3371/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_755 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3381 U$$3381/A _665_/Q VGND VGND VPWR VPWR U$$3381/X sky130_fd_sc_hd__xor2_1
XU$$3392 _600_/Q U$$3402/A2 _601_/Q U$$3402/B2 VGND VGND VPWR VPWR U$$3393/A sky130_fd_sc_hd__a22o_1
XFILLER_181_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_6_0 U$$19/X U$$152/X U$$285/X VGND VGND VPWR VPWR dadda_fa_6_7_0/A dadda_fa_6_6_0/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_90_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2680 U$$2680/A U$$2698/B VGND VGND VPWR VPWR U$$2680/X sky130_fd_sc_hd__xor2_1
XU$$2691 U$$4061/A1 U$$2733/A2 U$$3652/A1 U$$2733/B2 VGND VGND VPWR VPWR U$$2692/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_clk _535_/CLK VGND VGND VPWR VPWR _588_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1990 U$$757/A1 U$$2040/A2 U$$759/A1 U$$2040/B2 VGND VGND VPWR VPWR U$$1991/A sky130_fd_sc_hd__a22o_1
XFILLER_167_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_81_2 dadda_fa_4_81_2/A dadda_fa_4_81_2/B dadda_fa_4_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/CIN dadda_fa_5_81_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_190_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_74_1 dadda_fa_4_74_1/A dadda_fa_4_74_1/B dadda_fa_4_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/B dadda_fa_5_74_1/B sky130_fd_sc_hd__fa_1
XFILLER_116_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_51_0 dadda_fa_7_51_0/A dadda_fa_7_51_0/B dadda_fa_7_51_0/CIN VGND VGND
+ VPWR VPWR _476_/D _347_/D sky130_fd_sc_hd__fa_2
XFILLER_62_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_67_0 dadda_fa_4_67_0/A dadda_fa_4_67_0/B dadda_fa_4_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/A dadda_fa_5_67_1/A sky130_fd_sc_hd__fa_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput104 b[45] VGND VGND VPWR VPWR _597_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput115 b[55] VGND VGND VPWR VPWR _607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput126 b[7] VGND VGND VPWR VPWR _559_/D sky130_fd_sc_hd__clkbuf_1
XTAP_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput137 c[107] VGND VGND VPWR VPWR input137/X sky130_fd_sc_hd__clkbuf_2
XTAP_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput148 c[117] VGND VGND VPWR VPWR input148/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput159 c[127] VGND VGND VPWR VPWR input159/X sky130_fd_sc_hd__clkbuf_1
XTAP_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$631 final_adder.U$$9/SUM final_adder.U$$631/B VGND VGND VPWR VPWR
+ _177_/D sky130_fd_sc_hd__xor2_4
XTAP_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_640_ _648_/CLK _640_/D VGND VGND VPWR VPWR _640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$642 final_adder.U$$642/A final_adder.U$$642/B VGND VGND VPWR VPWR
+ _188_/D sky130_fd_sc_hd__xor2_4
XTAP_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$653 final_adder.U$$653/A final_adder.U$$653/B VGND VGND VPWR VPWR
+ _199_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$664 final_adder.U$$664/A final_adder.U$$664/B VGND VGND VPWR VPWR
+ _210_/D sky130_fd_sc_hd__xor2_2
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$503 U$$912/B1 U$$517/A2 U$$914/B1 U$$517/B2 VGND VGND VPWR VPWR U$$504/A sky130_fd_sc_hd__a22o_1
XFILLER_57_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$675 final_adder.U$$675/A final_adder.U$$675/B VGND VGND VPWR VPWR
+ _221_/D sky130_fd_sc_hd__xor2_1
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$514 U$$514/A U$$518/B VGND VGND VPWR VPWR U$$514/X sky130_fd_sc_hd__xor2_1
XFILLER_57_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$686 final_adder.U$$686/A final_adder.U$$686/B VGND VGND VPWR VPWR
+ _232_/D sky130_fd_sc_hd__xor2_1
XFILLER_186_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$525 U$$525/A1 U$$545/A2 U$$527/A1 U$$545/B2 VGND VGND VPWR VPWR U$$526/A sky130_fd_sc_hd__a22o_1
X_571_ _575_/CLK _571_/D VGND VGND VPWR VPWR _571_/Q sky130_fd_sc_hd__dfxtp_2
Xrepeater890 U$$62/B2 VGND VGND VPWR VPWR U$$68/B2 sky130_fd_sc_hd__buf_6
XFILLER_5_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$697 final_adder.U$$697/A final_adder.U$$697/B VGND VGND VPWR VPWR
+ _243_/D sky130_fd_sc_hd__xor2_2
XU$$536 U$$536/A U$$536/B VGND VGND VPWR VPWR U$$536/X sky130_fd_sc_hd__xor2_1
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$547 U$$547/A VGND VGND VPWR VPWR U$$547/Y sky130_fd_sc_hd__inv_1
XFILLER_147_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$558 U$$695/A1 U$$574/A2 U$$695/B1 U$$574/B2 VGND VGND VPWR VPWR U$$559/A sky130_fd_sc_hd__a22o_1
XFILLER_204_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$569 U$$569/A U$$665/B VGND VGND VPWR VPWR U$$569/X sky130_fd_sc_hd__xor2_1
XFILLER_32_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk _369_/CLK VGND VGND VPWR VPWR _520_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_201_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_444 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1403 U$$3916/B1 VGND VGND VPWR VPWR U$$80/B1 sky130_fd_sc_hd__buf_4
Xrepeater1414 U$$4053/A1 VGND VGND VPWR VPWR U$$628/A1 sky130_fd_sc_hd__buf_6
XFILLER_67_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1425 U$$4462/A1 VGND VGND VPWR VPWR U$$3503/A1 sky130_fd_sc_hd__clkbuf_8
Xrepeater1436 U$$4184/A1 VGND VGND VPWR VPWR U$$896/A1 sky130_fd_sc_hd__buf_6
XFILLER_153_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1447 _584_/Q VGND VGND VPWR VPWR U$$4317/B1 sky130_fd_sc_hd__clkbuf_8
Xrepeater1458 _583_/Q VGND VGND VPWR VPWR U$$4180/A1 sky130_fd_sc_hd__buf_6
Xrepeater1469 U$$3626/B1 VGND VGND VPWR VPWR U$$749/B1 sky130_fd_sc_hd__buf_8
XFILLER_137_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$5_1838 VGND VGND VPWR VPWR U$$5_1838/HI U$$5/A2 sky130_fd_sc_hd__conb_1
XFILLER_67_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1220 U$$2588/B1 U$$1224/A2 U$$948/A1 U$$1224/B2 VGND VGND VPWR VPWR U$$1221/A
+ sky130_fd_sc_hd__a22o_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1231 U$$1231/A U$$1232/A VGND VGND VPWR VPWR U$$1231/X sky130_fd_sc_hd__xor2_1
XFILLER_206_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1242 U$$1242/A U$$1296/B VGND VGND VPWR VPWR U$$1242/X sky130_fd_sc_hd__xor2_1
XU$$1253 U$$840/B1 U$$1291/A2 U$$568/B1 U$$1291/B2 VGND VGND VPWR VPWR U$$1254/A sky130_fd_sc_hd__a22o_1
XU$$1264 U$$1264/A U$$1292/B VGND VGND VPWR VPWR U$$1264/X sky130_fd_sc_hd__xor2_1
XU$$1275 U$$2508/A1 U$$1279/A2 U$$2508/B1 U$$1279/B2 VGND VGND VPWR VPWR U$$1276/A
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_42_clk _369_/CLK VGND VGND VPWR VPWR _510_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1286 U$$1286/A U$$1332/B VGND VGND VPWR VPWR U$$1286/X sky130_fd_sc_hd__xor2_1
XU$$1297 U$$749/A1 U$$1309/A2 U$$749/B1 U$$1309/B2 VGND VGND VPWR VPWR U$$1298/A sky130_fd_sc_hd__a22o_1
XFILLER_31_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_91_1 dadda_fa_5_91_1/A dadda_fa_5_91_1/B dadda_fa_5_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_92_0/B dadda_fa_7_91_0/A sky130_fd_sc_hd__fa_1
XFILLER_191_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_84_0 dadda_fa_5_84_0/A dadda_fa_5_84_0/B dadda_fa_5_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_85_0/A dadda_fa_6_84_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_76_7 U$$4282/X U$$4415/X input230/X VGND VGND VPWR VPWR dadda_fa_2_77_2/CIN
+ dadda_fa_2_76_5/CIN sky130_fd_sc_hd__fa_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_6 dadda_fa_1_69_6/A dadda_fa_1_69_6/B dadda_fa_1_69_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_2/B dadda_fa_2_69_5/B sky130_fd_sc_hd__fa_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_clk _479_/CLK VGND VGND VPWR VPWR _351_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_99_0 dadda_fa_7_99_0/A dadda_fa_7_99_0/B dadda_fa_7_99_0/CIN VGND VGND
+ VPWR VPWR _524_/D _395_/D sky130_fd_sc_hd__fa_1
XFILLER_139_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_786 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_47 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_100_2 dadda_fa_3_100_2/A dadda_fa_3_100_2/B dadda_fa_3_100_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_1/A dadda_fa_4_100_2/B sky130_fd_sc_hd__fa_1
XFILLER_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_803 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_64_5 U$$2130/X U$$2263/X U$$2396/X VGND VGND VPWR VPWR dadda_fa_1_65_7/A
+ dadda_fa_2_64_0/A sky130_fd_sc_hd__fa_2
XTAP_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_114_0 dadda_fa_6_114_0/A dadda_fa_6_114_0/B dadda_fa_6_114_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_115_0/B dadda_fa_7_114_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_40_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$300 U$$26/A1 U$$308/A2 U$$28/A1 U$$308/B2 VGND VGND VPWR VPWR U$$301/A sky130_fd_sc_hd__a22o_1
XFILLER_18_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$461 final_adder.U$$284/B final_adder.U$$678/B final_adder.U$$185/X
+ VGND VGND VPWR VPWR final_adder.U$$680/B sky130_fd_sc_hd__a21o_1
XTAP_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_623_ _623_/CLK _623_/D VGND VGND VPWR VPWR _623_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$311 U$$311/A U$$319/B VGND VGND VPWR VPWR U$$311/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$483 final_adder.U$$306/B final_adder.U$$722/B final_adder.U$$229/X
+ VGND VGND VPWR VPWR final_adder.U$$724/B sky130_fd_sc_hd__a21o_1
Xdadda_fa_3_34_3 dadda_fa_3_34_3/A dadda_fa_3_34_3/B dadda_fa_3_34_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_1/B dadda_fa_4_34_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$322 U$$733/A1 U$$334/A2 U$$733/B1 U$$334/B2 VGND VGND VPWR VPWR U$$323/A sky130_fd_sc_hd__a22o_1
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$333 U$$333/A U$$397/B VGND VGND VPWR VPWR U$$333/X sky130_fd_sc_hd__xor2_1
XFILLER_44_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$344 U$$344/A1 U$$350/A2 U$$72/A1 U$$350/B2 VGND VGND VPWR VPWR U$$345/A sky130_fd_sc_hd__a22o_1
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_27_2 input176/X dadda_fa_3_27_2/B dadda_fa_3_27_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_28_1/A dadda_fa_4_27_2/B sky130_fd_sc_hd__fa_1
XU$$355 U$$355/A U$$397/B VGND VGND VPWR VPWR U$$355/X sky130_fd_sc_hd__xor2_1
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_554_ _558_/CLK _554_/D VGND VGND VPWR VPWR _554_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$366 U$$912/B1 U$$392/A2 U$$368/A1 U$$392/B2 VGND VGND VPWR VPWR U$$367/A sky130_fd_sc_hd__a22o_1
XU$$377 U$$377/A U$$383/B VGND VGND VPWR VPWR U$$377/X sky130_fd_sc_hd__xor2_1
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$388 U$$525/A1 U$$392/A2 U$$527/A1 U$$392/B2 VGND VGND VPWR VPWR U$$389/A sky130_fd_sc_hd__a22o_1
XU$$399 U$$399/A U$$411/A VGND VGND VPWR VPWR U$$399/X sky130_fd_sc_hd__xor2_1
Xclkbuf_2_3_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_3_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_485_ _485_/CLK _485_/D VGND VGND VPWR VPWR _485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_clk _432_/CLK VGND VGND VPWR VPWR _189_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1200 U$$954/A1 VGND VGND VPWR VPWR U$$817/A1 sky130_fd_sc_hd__buf_6
XFILLER_172_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1211 U$$952/A1 VGND VGND VPWR VPWR U$$3418/A1 sky130_fd_sc_hd__buf_6
Xrepeater1222 U$$3005/A1 VGND VGND VPWR VPWR U$$2318/B1 sky130_fd_sc_hd__buf_6
Xrepeater1233 U$$2314/B1 VGND VGND VPWR VPWR U$$944/B1 sky130_fd_sc_hd__buf_4
Xrepeater1244 U$$4506/A1 VGND VGND VPWR VPWR U$$4369/A1 sky130_fd_sc_hd__buf_4
Xrepeater1255 _608_/Q VGND VGND VPWR VPWR U$$3269/B1 sky130_fd_sc_hd__buf_4
XFILLER_99_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1266 U$$2171/A1 VGND VGND VPWR VPWR U$$527/A1 sky130_fd_sc_hd__buf_8
XFILLER_4_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1277 U$$4498/A1 VGND VGND VPWR VPWR U$$4224/A1 sky130_fd_sc_hd__buf_6
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1288 U$$3674/A1 VGND VGND VPWR VPWR U$$2715/A1 sky130_fd_sc_hd__buf_4
XFILLER_10_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1299 _602_/Q VGND VGND VPWR VPWR U$$3122/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_79_5 dadda_fa_2_79_5/A dadda_fa_2_79_5/B dadda_fa_2_79_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_2/A dadda_fa_4_79_0/A sky130_fd_sc_hd__fa_2
XFILLER_84_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_30_4 U$$1663/X U$$1796/X VGND VGND VPWR VPWR dadda_fa_3_31_2/B dadda_fa_4_30_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_7_0_0 U$$7/X U$$9/B VGND VGND VPWR VPWR _425_/D _296_/D sky130_fd_sc_hd__ha_1
XFILLER_36_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1050 U$$1050/A U$$1090/B VGND VGND VPWR VPWR U$$1050/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_15_clk _616_/CLK VGND VGND VPWR VPWR _487_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_211_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1061 U$$2705/A1 U$$1065/A2 U$$926/A1 U$$1065/B2 VGND VGND VPWR VPWR U$$1062/A
+ sky130_fd_sc_hd__a22o_1
XU$$1072 U$$1072/A U$$1078/B VGND VGND VPWR VPWR U$$1072/X sky130_fd_sc_hd__xor2_1
XFILLER_32_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1083 U$$946/A1 U$$1093/A2 U$$946/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1084/A sky130_fd_sc_hd__a22o_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1094 U$$1094/A U$$1095/A VGND VGND VPWR VPWR U$$1094/X sky130_fd_sc_hd__xor2_1
XFILLER_148_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_82_7 U$$4028/X U$$4161/X VGND VGND VPWR VPWR dadda_fa_2_83_3/CIN dadda_fa_3_82_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_109_1 dadda_fa_5_109_1/A dadda_fa_5_109_1/B dadda_fa_5_109_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_110_0/B dadda_fa_7_109_0/A sky130_fd_sc_hd__fa_1
XFILLER_117_543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_81_5 U$$3228/X U$$3361/X U$$3494/X VGND VGND VPWR VPWR dadda_fa_2_82_2/CIN
+ dadda_fa_2_81_5/B sky130_fd_sc_hd__fa_1
XFILLER_63_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_74_4 U$$3347/X U$$3480/X U$$3613/X VGND VGND VPWR VPWR dadda_fa_2_75_1/CIN
+ dadda_fa_2_74_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_67_3 U$$3732/X U$$3865/X U$$3998/X VGND VGND VPWR VPWR dadda_fa_2_68_1/B
+ dadda_fa_2_67_4/B sky130_fd_sc_hd__fa_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_44_2 dadda_fa_4_44_2/A dadda_fa_4_44_2/B dadda_fa_4_44_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/CIN dadda_fa_5_44_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_37_1 dadda_fa_4_37_1/A dadda_fa_4_37_1/B dadda_fa_4_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/B dadda_fa_5_37_1/B sky130_fd_sc_hd__fa_1
XFILLER_160_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_14_0 dadda_fa_7_14_0/A dadda_fa_7_14_0/B dadda_fa_7_14_0/CIN VGND VGND
+ VPWR VPWR _439_/D _310_/D sky130_fd_sc_hd__fa_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_270_ _520_/CLK _270_/D VGND VGND VPWR VPWR _270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_332 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_62_2 U$$929/X U$$1062/X U$$1195/X VGND VGND VPWR VPWR dadda_fa_1_63_6/A
+ dadda_fa_1_62_8/A sky130_fd_sc_hd__fa_1
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3903 U$$3903/A U$$3949/B VGND VGND VPWR VPWR U$$3903/X sky130_fd_sc_hd__xor2_1
XFILLER_76_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3914 U$$4462/A1 U$$3916/A2 U$$4464/A1 U$$3916/B2 VGND VGND VPWR VPWR U$$3915/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3925 U$$3925/A U$$3935/B VGND VGND VPWR VPWR U$$3925/X sky130_fd_sc_hd__xor2_1
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_338 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3936 U$$4208/B1 U$$3840/X U$$4075/A1 U$$3841/X VGND VGND VPWR VPWR U$$3937/A sky130_fd_sc_hd__a22o_1
XU$$3947 U$$3947/A U$$3973/A VGND VGND VPWR VPWR U$$3947/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_32_0 U$$2263/B input182/X dadda_fa_3_32_0/CIN VGND VGND VPWR VPWR dadda_fa_4_33_0/B
+ dadda_fa_4_32_1/CIN sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$280 final_adder.U$$280/A final_adder.U$$280/B VGND VGND VPWR VPWR
+ final_adder.U$$332/B sky130_fd_sc_hd__and2_1
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3958 U$$4369/A1 U$$3958/A2 U$$4369/B1 U$$3958/B2 VGND VGND VPWR VPWR U$$3959/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_606_ _613_/CLK _606_/D VGND VGND VPWR VPWR _606_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3969 U$$3969/A U$$3973/A VGND VGND VPWR VPWR U$$3969/X sky130_fd_sc_hd__xor2_1
XU$$130 U$$676/B1 U$$4/X U$$406/A1 U$$5/X VGND VGND VPWR VPWR U$$131/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$291 final_adder.U$$290/A final_adder.U$$197/X final_adder.U$$199/X
+ VGND VGND VPWR VPWR final_adder.U$$291/X sky130_fd_sc_hd__a21o_1
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$141 U$$139/Y _618_/Q U$$2/A U$$140/X U$$137/Y VGND VGND VPWR VPWR U$$141/X sky130_fd_sc_hd__a32o_1
XFILLER_33_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$152 U$$152/A U$$180/B VGND VGND VPWR VPWR U$$152/X sky130_fd_sc_hd__xor2_1
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$163 U$$26/A1 U$$175/A2 U$$28/A1 U$$175/B2 VGND VGND VPWR VPWR U$$164/A sky130_fd_sc_hd__a22o_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$174 U$$174/A U$$196/B VGND VGND VPWR VPWR U$$174/X sky130_fd_sc_hd__xor2_1
X_537_ _538_/CLK _537_/D VGND VGND VPWR VPWR _537_/Q sky130_fd_sc_hd__dfxtp_1
XU$$185 U$$733/A1 U$$219/A2 U$$50/A1 U$$219/B2 VGND VGND VPWR VPWR U$$186/A sky130_fd_sc_hd__a22o_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$196 U$$196/A U$$196/B VGND VGND VPWR VPWR U$$196/X sky130_fd_sc_hd__xor2_1
XFILLER_60_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_468_ _471_/CLK _468_/D VGND VGND VPWR VPWR _468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_399_ _526_/CLK _399_/D VGND VGND VPWR VPWR _399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_91_4 dadda_fa_2_91_4/A dadda_fa_2_91_4/B dadda_fa_2_91_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_92_1/CIN dadda_fa_3_91_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_57_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1030 U$$2465/A VGND VGND VPWR VPWR U$$2462/B sky130_fd_sc_hd__buf_6
Xrepeater1041 U$$2303/B VGND VGND VPWR VPWR U$$2299/B sky130_fd_sc_hd__buf_6
XFILLER_99_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1052 U$$2174/B VGND VGND VPWR VPWR U$$2170/B sky130_fd_sc_hd__buf_6
XFILLER_86_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1063 _645_/Q VGND VGND VPWR VPWR U$$2043/B sky130_fd_sc_hd__buf_8
Xdadda_fa_2_84_3 dadda_fa_2_84_3/A dadda_fa_2_84_3/B dadda_fa_2_84_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/B dadda_fa_3_84_3/B sky130_fd_sc_hd__fa_1
XFILLER_153_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1074 U$$1737/B VGND VGND VPWR VPWR U$$1687/B sky130_fd_sc_hd__buf_6
Xrepeater1085 U$$1642/B VGND VGND VPWR VPWR U$$1598/B sky130_fd_sc_hd__buf_6
Xrepeater1096 U$$1479/B VGND VGND VPWR VPWR U$$1429/B sky130_fd_sc_hd__buf_12
Xdadda_fa_2_77_2 dadda_fa_2_77_2/A dadda_fa_2_77_2/B dadda_fa_2_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/A dadda_fa_3_77_3/A sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_4_clk _442_/CLK VGND VGND VPWR VPWR _469_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_5_54_1 dadda_fa_5_54_1/A dadda_fa_5_54_1/B dadda_fa_5_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_55_0/B dadda_fa_7_54_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_47_0 dadda_fa_5_47_0/A dadda_fa_5_47_0/B dadda_fa_5_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_48_0/A dadda_fa_6_47_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_210_1109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_100_1 U$$2867/X U$$3000/X U$$3133/X VGND VGND VPWR VPWR dadda_fa_3_101_1/CIN
+ dadda_fa_3_100_3/A sky130_fd_sc_hd__fa_1
XFILLER_36_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_121_0 U$$4372/X U$$4505/X input153/X VGND VGND VPWR VPWR dadda_fa_6_122_0/A
+ dadda_fa_6_121_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_72_1 U$$2412/X U$$2545/X U$$2678/X VGND VGND VPWR VPWR dadda_fa_2_73_0/CIN
+ dadda_fa_2_72_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_931 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_590 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_65_0 U$$2531/X U$$2664/X U$$2797/X VGND VGND VPWR VPWR dadda_fa_2_66_0/B
+ dadda_fa_2_65_3/B sky130_fd_sc_hd__fa_1
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_614 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2509 U$$2509/A U$$2551/B VGND VGND VPWR VPWR U$$2509/X sky130_fd_sc_hd__xor2_1
XFILLER_62_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1808 U$$1808/A U$$1844/B VGND VGND VPWR VPWR U$$1808/X sky130_fd_sc_hd__xor2_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1819 U$$38/A1 U$$1859/A2 U$$40/A1 U$$1859/B2 VGND VGND VPWR VPWR U$$1820/A sky130_fd_sc_hd__a22o_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ _451_/CLK _322_/D VGND VGND VPWR VPWR _322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_920 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_253_ _253_/CLK _253_/D VGND VGND VPWR VPWR _253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_986 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_184_ _189_/CLK _184_/D VGND VGND VPWR VPWR _184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_94_2 dadda_fa_3_94_2/A dadda_fa_3_94_2/B dadda_fa_3_94_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_1/A dadda_fa_4_94_2/B sky130_fd_sc_hd__fa_1
XFILLER_171_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_87_1 dadda_fa_3_87_1/A dadda_fa_3_87_1/B dadda_fa_3_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_0/CIN dadda_fa_4_87_2/A sky130_fd_sc_hd__fa_1
XFILLER_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_64_0 dadda_fa_6_64_0/A dadda_fa_6_64_0/B dadda_fa_6_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_65_0/B dadda_fa_7_64_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_9_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater708 U$$3968/B2 VGND VGND VPWR VPWR U$$3958/B2 sky130_fd_sc_hd__buf_6
XFILLER_81_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater719 U$$3674/B2 VGND VGND VPWR VPWR U$$3628/B2 sky130_fd_sc_hd__buf_4
XU$$4401 U$$4401/A U$$4401/B VGND VGND VPWR VPWR U$$4401/X sky130_fd_sc_hd__xor2_1
XU$$4412 _562_/Q U$$4388/X _563_/Q U$$4430/B2 VGND VGND VPWR VPWR U$$4413/A sky130_fd_sc_hd__a22o_1
XU$$4423 U$$4423/A U$$4423/B VGND VGND VPWR VPWR U$$4423/X sky130_fd_sc_hd__xor2_1
XFILLER_78_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4434 U$$4434/A1 U$$4388/X _574_/Q U$$4438/B2 VGND VGND VPWR VPWR U$$4435/A sky130_fd_sc_hd__a22o_1
XFILLER_77_474 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4431_1794 VGND VGND VPWR VPWR U$$4431_1794/HI U$$4431/B sky130_fd_sc_hd__conb_1
XFILLER_49_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3700 _670_/Q VGND VGND VPWR VPWR U$$3702/B sky130_fd_sc_hd__inv_1
XFILLER_92_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4445 U$$4445/A U$$4445/B VGND VGND VPWR VPWR U$$4445/X sky130_fd_sc_hd__xor2_1
XU$$4456 _584_/Q U$$4388/X U$$4456/B1 U$$4468/B2 VGND VGND VPWR VPWR U$$4457/A sky130_fd_sc_hd__a22o_1
XU$$3711 _554_/Q U$$3743/A2 U$$3713/A1 U$$3743/B2 VGND VGND VPWR VPWR U$$3712/A sky130_fd_sc_hd__a22o_1
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_116_1 U$$4229/X U$$4362/X U$$4495/X VGND VGND VPWR VPWR dadda_fa_5_117_0/B
+ dadda_fa_5_116_1/B sky130_fd_sc_hd__fa_1
XFILLER_37_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3722 U$$3722/A U$$3740/B VGND VGND VPWR VPWR U$$3722/X sky130_fd_sc_hd__xor2_1
XFILLER_65_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4467 U$$4467/A U$$4467/B VGND VGND VPWR VPWR U$$4467/X sky130_fd_sc_hd__xor2_1
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3733 _565_/Q U$$3769/A2 U$$3735/A1 U$$3769/B2 VGND VGND VPWR VPWR U$$3734/A sky130_fd_sc_hd__a22o_1
XFILLER_53_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4478 U$$4478/A1 U$$4388/X U$$4480/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4479/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3744 U$$3744/A U$$3764/B VGND VGND VPWR VPWR U$$3744/X sky130_fd_sc_hd__xor2_1
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4489 U$$4489/A U$$4489/B VGND VGND VPWR VPWR U$$4489/X sky130_fd_sc_hd__xor2_1
XFILLER_93_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_7__f_clk clkbuf_2_3_0_clk/X VGND VGND VPWR VPWR _535_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$3755 _576_/Q U$$3785/A2 _577_/Q U$$3785/B2 VGND VGND VPWR VPWR U$$3756/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_109_0 dadda_fa_4_109_0/A dadda_fa_4_109_0/B dadda_fa_4_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/A dadda_fa_5_109_1/A sky130_fd_sc_hd__fa_1
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3766 U$$3766/A _671_/Q VGND VGND VPWR VPWR U$$3766/X sky130_fd_sc_hd__xor2_1
XU$$3777 U$$4462/A1 U$$3777/A2 U$$4464/A1 U$$3777/B2 VGND VGND VPWR VPWR U$$3778/A
+ sky130_fd_sc_hd__a22o_1
XU$$3788 U$$3788/A U$$3804/B VGND VGND VPWR VPWR U$$3788/X sky130_fd_sc_hd__xor2_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4507_1832 VGND VGND VPWR VPWR U$$4507_1832/HI U$$4507/B sky130_fd_sc_hd__conb_1
XU$$3799 U$$3934/B1 U$$3805/A2 U$$3799/B1 U$$3805/B2 VGND VGND VPWR VPWR U$$3800/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_370 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_381 U$$429/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_392 U$$1922/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_82_0 U$$4294/X U$$4427/X input237/X VGND VGND VPWR VPWR dadda_fa_3_83_0/B
+ dadda_fa_3_82_2/B sky130_fd_sc_hd__fa_1
XFILLER_142_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_51_6 U$$2503/X U$$2636/X U$$2769/X VGND VGND VPWR VPWR dadda_fa_2_52_2/B
+ dadda_fa_2_51_5/B sky130_fd_sc_hd__fa_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_3_0 input190/X dadda_fa_7_3_0/B dadda_ha_6_3_0/SUM VGND VGND VPWR VPWR
+ _428_/D _299_/D sky130_fd_sc_hd__fa_1
XFILLER_37_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_582 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_755 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_81_0 dadda_fa_7_81_0/A dadda_fa_7_81_0/B dadda_fa_7_81_0/CIN VGND VGND
+ VPWR VPWR _506_/D _377_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_97_0 dadda_fa_4_97_0/A dadda_fa_4_97_0/B dadda_fa_4_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/A dadda_fa_5_97_1/A sky130_fd_sc_hd__fa_1
XFILLER_152_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_271 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3007 U$$3281/A1 U$$2881/X U$$3283/A1 U$$2882/X VGND VGND VPWR VPWR U$$3008/A sky130_fd_sc_hd__a22o_1
XU$$3018 U$$3016/Y _660_/Q U$$3014/A U$$3017/X U$$3014/Y VGND VGND VPWR VPWR U$$3018/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3029 U$$3029/A U$$3077/B VGND VGND VPWR VPWR U$$3029/X sky130_fd_sc_hd__xor2_1
XU$$2306 U$$4224/A1 U$$2196/X U$$4361/B1 U$$2197/X VGND VGND VPWR VPWR U$$2307/A sky130_fd_sc_hd__a22o_1
XU$$2317 U$$2317/A U$$2321/B VGND VGND VPWR VPWR U$$2317/X sky130_fd_sc_hd__xor2_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2328 U$$2328/A VGND VGND VPWR VPWR U$$2328/Y sky130_fd_sc_hd__inv_1
XFILLER_90_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2339 U$$2611/B1 U$$2367/A2 U$$2478/A1 U$$2367/B2 VGND VGND VPWR VPWR U$$2340/A
+ sky130_fd_sc_hd__a22o_1
XU$$1605 U$$3112/A1 U$$1607/A2 U$$922/A1 U$$1607/B2 VGND VGND VPWR VPWR U$$1606/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1616 U$$1616/A U$$1636/B VGND VGND VPWR VPWR U$$1616/X sky130_fd_sc_hd__xor2_1
XFILLER_27_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1627 U$$2721/B1 U$$1627/A2 U$$2586/B1 U$$1627/B2 VGND VGND VPWR VPWR U$$1628/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1638 U$$1638/A _639_/Q VGND VGND VPWR VPWR U$$1638/X sky130_fd_sc_hd__xor2_1
XFILLER_203_634 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1649 U$$1647/B _639_/Q _640_/Q U$$1644/Y VGND VGND VPWR VPWR U$$1649/X sky130_fd_sc_hd__a22o_2
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_396 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_305_ _435_/CLK _305_/D VGND VGND VPWR VPWR _305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_236_ _503_/CLK _236_/D VGND VGND VPWR VPWR _236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_61_5 dadda_fa_2_61_5/A dadda_fa_2_61_5/B dadda_fa_2_61_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_2/A dadda_fa_4_61_0/A sky130_fd_sc_hd__fa_2
Xrepeater505 U$$3110/A2 VGND VGND VPWR VPWR U$$3082/A2 sky130_fd_sc_hd__buf_8
Xrepeater516 U$$3005/A2 VGND VGND VPWR VPWR U$$2981/A2 sky130_fd_sc_hd__buf_12
Xrepeater527 U$$2812/A2 VGND VGND VPWR VPWR U$$2814/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_54_4 dadda_fa_2_54_4/A dadda_fa_2_54_4/B dadda_fa_2_54_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/CIN dadda_fa_3_54_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_ha_2_108_0_1875 VGND VGND VPWR VPWR dadda_ha_2_108_0/A dadda_ha_2_108_0_1875/LO
+ sky130_fd_sc_hd__conb_1
Xrepeater538 U$$2707/A2 VGND VGND VPWR VPWR U$$2705/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4220 U$$4355/B1 U$$4238/A2 U$$4222/A1 U$$4238/B2 VGND VGND VPWR VPWR U$$4221/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater549 U$$2580/A2 VGND VGND VPWR VPWR U$$2588/A2 sky130_fd_sc_hd__buf_6
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4231 U$$4231/A U$$4239/B VGND VGND VPWR VPWR U$$4231/X sky130_fd_sc_hd__xor2_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4242 U$$4516/A1 U$$4244/A2 U$$4516/B1 U$$4244/B2 VGND VGND VPWR VPWR U$$4243/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4253 U$$4253/A1 U$$4297/A2 U$$4392/A1 U$$4297/B2 VGND VGND VPWR VPWR U$$4254/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_47_3 dadda_fa_2_47_3/A dadda_fa_2_47_3/B dadda_fa_2_47_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/B dadda_fa_3_47_3/B sky130_fd_sc_hd__fa_1
XU$$4264 U$$4264/A U$$4348/B VGND VGND VPWR VPWR U$$4264/X sky130_fd_sc_hd__xor2_1
XU$$3530 U$$3530/A U$$3538/B VGND VGND VPWR VPWR U$$3530/X sky130_fd_sc_hd__xor2_1
XU$$4275 _562_/Q U$$4311/A2 _563_/Q U$$4311/B2 VGND VGND VPWR VPWR U$$4276/A sky130_fd_sc_hd__a22o_1
XU$$4286 U$$4286/A U$$4322/B VGND VGND VPWR VPWR U$$4286/X sky130_fd_sc_hd__xor2_1
XFILLER_53_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3541 U$$4087/B1 U$$3555/A2 U$$3952/B1 U$$3555/B2 VGND VGND VPWR VPWR U$$3542/A
+ sky130_fd_sc_hd__a22o_1
XU$$3552 U$$3552/A U$$3556/B VGND VGND VPWR VPWR U$$3552/X sky130_fd_sc_hd__xor2_1
XU$$4297 _573_/Q U$$4297/A2 _574_/Q U$$4297/B2 VGND VGND VPWR VPWR U$$4298/A sky130_fd_sc_hd__a22o_1
XU$$3563 _668_/Q VGND VGND VPWR VPWR U$$3565/B sky130_fd_sc_hd__inv_1
XFILLER_20_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3574 _554_/Q U$$3612/A2 U$$3713/A1 U$$3612/B2 VGND VGND VPWR VPWR U$$3575/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_17_1 dadda_fa_5_17_1/A dadda_fa_5_17_1/B dadda_fa_5_17_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_18_0/B dadda_fa_7_17_0/A sky130_fd_sc_hd__fa_1
XU$$2840 U$$4208/B1 U$$2874/A2 U$$4075/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2841/A
+ sky130_fd_sc_hd__a22o_1
XU$$3585 U$$3585/A U$$3609/B VGND VGND VPWR VPWR U$$3585/X sky130_fd_sc_hd__xor2_1
XU$$2851 U$$2851/A _657_/Q VGND VGND VPWR VPWR U$$2851/X sky130_fd_sc_hd__xor2_1
XU$$3596 _565_/Q U$$3636/A2 U$$3735/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3597/A sky130_fd_sc_hd__a22o_1
XU$$2862 _609_/Q U$$2866/A2 U$$2999/B1 U$$2866/B2 VGND VGND VPWR VPWR U$$2863/A sky130_fd_sc_hd__a22o_1
XFILLER_45_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2873 U$$2873/A U$$2875/B VGND VGND VPWR VPWR U$$2873/X sky130_fd_sc_hd__xor2_1
XU$$2884 U$$2884/A U$$2928/B VGND VGND VPWR VPWR U$$2884/X sky130_fd_sc_hd__xor2_1
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2895 U$$2895/A1 U$$2943/A2 U$$3717/B1 U$$2943/B2 VGND VGND VPWR VPWR U$$2896/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1069 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_4_120_1 U$$4237/X U$$4370/X VGND VGND VPWR VPWR dadda_fa_5_121_1/B dadda_ha_4_120_1/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_143_972 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_43_4 U$$1689/X U$$1822/X VGND VGND VPWR VPWR dadda_fa_2_44_4/A dadda_fa_3_43_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_25_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_4_13_2 U$$831/X input161/X VGND VGND VPWR VPWR dadda_fa_5_14_0/CIN dadda_ha_4_13_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_99_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$707 U$$707/A1 U$$725/A2 U$$22/B1 U$$725/B2 VGND VGND VPWR VPWR U$$708/A sky130_fd_sc_hd__a22o_1
XU$$718 U$$718/A U$$760/B VGND VGND VPWR VPWR U$$718/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_42_2 U$$889/X U$$1022/X U$$1155/X VGND VGND VPWR VPWR dadda_fa_2_43_3/CIN
+ dadda_fa_2_42_5/B sky130_fd_sc_hd__fa_1
XU$$729 U$$42/B1 U$$795/A2 U$$729/B1 U$$795/B2 VGND VGND VPWR VPWR U$$730/A sky130_fd_sc_hd__a22o_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_12_0 U$$31/X U$$164/X U$$297/X VGND VGND VPWR VPWR dadda_fa_5_13_0/A dadda_fa_5_12_1/A
+ sky130_fd_sc_hd__fa_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1607 U$$4140/B1 VGND VGND VPWR VPWR U$$3320/A1 sky130_fd_sc_hd__buf_6
XFILLER_193_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1618 _563_/Q VGND VGND VPWR VPWR U$$3042/B1 sky130_fd_sc_hd__buf_6
XFILLER_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1629 U$$985/A1 VGND VGND VPWR VPWR U$$26/A1 sky130_fd_sc_hd__buf_4
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_64_3 dadda_fa_3_64_3/A dadda_fa_3_64_3/B dadda_fa_3_64_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_1/B dadda_fa_4_64_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_57_2 dadda_fa_3_57_2/A dadda_fa_3_57_2/B dadda_fa_3_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_1/A dadda_fa_4_57_2/B sky130_fd_sc_hd__fa_1
XFILLER_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_27_0 dadda_fa_6_27_0/A dadda_fa_6_27_0/B dadda_fa_6_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_28_0/B dadda_fa_7_27_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2103 U$$2375/B1 U$$2109/A2 U$$3884/B1 U$$2109/B2 VGND VGND VPWR VPWR U$$2104/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2114 U$$2114/A U$$2170/B VGND VGND VPWR VPWR U$$2114/X sky130_fd_sc_hd__xor2_1
XU$$2125 U$$890/B1 U$$2135/A2 U$$757/A1 U$$2135/B2 VGND VGND VPWR VPWR U$$2126/A sky130_fd_sc_hd__a22o_1
XU$$2136 U$$2136/A U$$2136/B VGND VGND VPWR VPWR U$$2136/X sky130_fd_sc_hd__xor2_1
XU$$1402 U$$715/B1 U$$1442/A2 U$$582/A1 U$$1442/B2 VGND VGND VPWR VPWR U$$1403/A sky130_fd_sc_hd__a22o_1
XU$$2147 U$$914/A1 U$$2169/A2 U$$916/A1 U$$2169/B2 VGND VGND VPWR VPWR U$$2148/A sky130_fd_sc_hd__a22o_1
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2158 U$$2158/A U$$2191/A VGND VGND VPWR VPWR U$$2158/X sky130_fd_sc_hd__xor2_1
XU$$1413 U$$1413/A U$$1429/B VGND VGND VPWR VPWR U$$1413/X sky130_fd_sc_hd__xor2_1
XFILLER_62_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1424 U$$54/A1 U$$1424/A2 U$$56/A1 U$$1424/B2 VGND VGND VPWR VPWR U$$1425/A sky130_fd_sc_hd__a22o_1
XFILLER_16_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2169 U$$525/A1 U$$2169/A2 U$$2171/A1 U$$2169/B2 VGND VGND VPWR VPWR U$$2170/A
+ sky130_fd_sc_hd__a22o_1
XU$$1435 U$$1435/A U$$1443/B VGND VGND VPWR VPWR U$$1435/X sky130_fd_sc_hd__xor2_1
XFILLER_31_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1446 U$$76/A1 U$$1486/A2 U$$3229/A1 U$$1486/B2 VGND VGND VPWR VPWR U$$1447/A sky130_fd_sc_hd__a22o_1
XFILLER_163_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1457 U$$1457/A U$$1459/B VGND VGND VPWR VPWR U$$1457/X sky130_fd_sc_hd__xor2_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1468 U$$2838/A1 U$$1474/A2 U$$2838/B1 U$$1474/B2 VGND VGND VPWR VPWR U$$1469/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1479 U$$1479/A U$$1479/B VGND VGND VPWR VPWR U$$1479/X sky130_fd_sc_hd__xor2_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_219_ _225_/CLK _219_/D VGND VGND VPWR VPWR _219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_983 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$109 _533_/Q _405_/Q VGND VGND VPWR VPWR final_adder.U$$237/B1 final_adder.U$$731/A
+ sky130_fd_sc_hd__ha_2
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_52_1 dadda_fa_2_52_1/A dadda_fa_2_52_1/B dadda_fa_2_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_0/CIN dadda_fa_3_52_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_731 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4050 U$$4050/A U$$4058/B VGND VGND VPWR VPWR U$$4050/X sky130_fd_sc_hd__xor2_1
XFILLER_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4061 U$$4061/A1 U$$4061/A2 _593_/Q U$$4061/B2 VGND VGND VPWR VPWR U$$4062/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_45_0 U$$2358/X U$$2491/X U$$2624/X VGND VGND VPWR VPWR dadda_fa_3_46_0/B
+ dadda_fa_3_45_2/B sky130_fd_sc_hd__fa_1
XFILLER_66_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4072 U$$4072/A U$$4072/B VGND VGND VPWR VPWR U$$4072/X sky130_fd_sc_hd__xor2_1
XU$$4083 U$$4355/B1 U$$4107/A2 U$$4222/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4084/A
+ sky130_fd_sc_hd__a22o_1
XU$$4094 U$$4094/A U$$4096/B VGND VGND VPWR VPWR U$$4094/X sky130_fd_sc_hd__xor2_1
XU$$3360 U$$4317/B1 U$$3378/A2 U$$3362/A1 U$$3378/B2 VGND VGND VPWR VPWR U$$3361/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3371 U$$3371/A U$$3424/A VGND VGND VPWR VPWR U$$3371/X sky130_fd_sc_hd__xor2_1
XFILLER_198_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3382 U$$3791/B1 U$$3404/A2 U$$3658/A1 U$$3404/B2 VGND VGND VPWR VPWR U$$3383/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3393 U$$3393/A U$$3397/B VGND VGND VPWR VPWR U$$3393/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2670 U$$2670/A U$$2706/B VGND VGND VPWR VPWR U$$2670/X sky130_fd_sc_hd__xor2_1
XU$$2681 U$$3229/A1 U$$2697/A2 U$$2957/A1 U$$2697/B2 VGND VGND VPWR VPWR U$$2682/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2692 U$$2692/A U$$2734/B VGND VGND VPWR VPWR U$$2692/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1980 U$$3213/A1 U$$2028/A2 U$$3352/A1 U$$2028/B2 VGND VGND VPWR VPWR U$$1981/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1991 U$$1991/A U$$2043/B VGND VGND VPWR VPWR U$$1991/X sky130_fd_sc_hd__xor2_1
XFILLER_194_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_74_2 dadda_fa_4_74_2/A dadda_fa_4_74_2/B dadda_fa_4_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/CIN dadda_fa_5_74_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_67_1 dadda_fa_4_67_1/A dadda_fa_4_67_1/B dadda_fa_4_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/B dadda_fa_5_67_1/B sky130_fd_sc_hd__fa_1
Xinput105 b[46] VGND VGND VPWR VPWR _598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput116 b[56] VGND VGND VPWR VPWR _608_/D sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_7_44_0 dadda_fa_7_44_0/A dadda_fa_7_44_0/B dadda_fa_7_44_0/CIN VGND VGND
+ VPWR VPWR _469_/D _340_/D sky130_fd_sc_hd__fa_1
XFILLER_76_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput127 b[8] VGND VGND VPWR VPWR _560_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_34_0 U$$75/X U$$208/X VGND VGND VPWR VPWR dadda_fa_2_35_5/CIN dadda_fa_3_34_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_9_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput138 c[108] VGND VGND VPWR VPWR input138/X sky130_fd_sc_hd__clkbuf_2
XTAP_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput149 c[118] VGND VGND VPWR VPWR input149/X sky130_fd_sc_hd__clkbuf_1
XTAP_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$621 final_adder.U$$748/A final_adder.U$$748/B final_adder.U$$621/B1
+ VGND VGND VPWR VPWR final_adder.U$$749/B sky130_fd_sc_hd__a21o_1
XTAP_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$632 final_adder.U$$632/A final_adder.U$$632/B VGND VGND VPWR VPWR
+ _178_/D sky130_fd_sc_hd__xor2_4
XFILLER_116_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$643 final_adder.U$$643/A final_adder.U$$643/B VGND VGND VPWR VPWR
+ _189_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$654 final_adder.U$$654/A final_adder.U$$654/B VGND VGND VPWR VPWR
+ _200_/D sky130_fd_sc_hd__xor2_1
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1041 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$665 final_adder.U$$665/A final_adder.U$$665/B VGND VGND VPWR VPWR
+ _211_/D sky130_fd_sc_hd__xor2_2
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$504 U$$504/A U$$518/B VGND VGND VPWR VPWR U$$504/X sky130_fd_sc_hd__xor2_1
XFILLER_17_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$676 final_adder.U$$676/A final_adder.U$$676/B VGND VGND VPWR VPWR
+ _222_/D sky130_fd_sc_hd__xor2_1
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$515 U$$650/B1 U$$517/A2 U$$515/B1 U$$517/B2 VGND VGND VPWR VPWR U$$516/A sky130_fd_sc_hd__a22o_1
X_570_ _572_/CLK _570_/D VGND VGND VPWR VPWR _570_/Q sky130_fd_sc_hd__dfxtp_4
Xrepeater880 U$$1190/B2 VGND VGND VPWR VPWR U$$1150/B2 sky130_fd_sc_hd__buf_6
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$526 U$$526/A U$$547/A VGND VGND VPWR VPWR U$$526/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$687 final_adder.U$$687/A final_adder.U$$687/B VGND VGND VPWR VPWR
+ _233_/D sky130_fd_sc_hd__xor2_4
Xrepeater891 U$$98/B2 VGND VGND VPWR VPWR U$$118/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$698 final_adder.U$$698/A final_adder.U$$698/B VGND VGND VPWR VPWR
+ _244_/D sky130_fd_sc_hd__xor2_1
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$537 U$$674/A1 U$$415/X U$$676/A1 U$$416/X VGND VGND VPWR VPWR U$$538/A sky130_fd_sc_hd__a22o_1
XFILLER_45_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$548 _623_/Q VGND VGND VPWR VPWR U$$548/Y sky130_fd_sc_hd__inv_1
XFILLER_205_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$559 U$$559/A U$$589/B VGND VGND VPWR VPWR U$$559/X sky130_fd_sc_hd__xor2_1
XFILLER_204_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1083 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1404 U$$82/A1 VGND VGND VPWR VPWR U$$493/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1415 U$$4053/A1 VGND VGND VPWR VPWR U$$2957/A1 sky130_fd_sc_hd__buf_8
XFILLER_197_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1426 _587_/Q VGND VGND VPWR VPWR U$$4462/A1 sky130_fd_sc_hd__buf_4
Xrepeater1437 U$$3362/A1 VGND VGND VPWR VPWR U$$759/A1 sky130_fd_sc_hd__buf_4
XFILLER_193_1026 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1448 U$$3769/B1 VGND VGND VPWR VPWR U$$757/A1 sky130_fd_sc_hd__buf_4
Xrepeater1459 U$$68/A1 VGND VGND VPWR VPWR U$$614/B1 sky130_fd_sc_hd__buf_6
XFILLER_158_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_75 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_62_0 dadda_fa_3_62_0/A dadda_fa_3_62_0/B dadda_fa_3_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_0/B dadda_fa_4_62_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_252 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_583 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_4_9_0 U$$25/X U$$158/X VGND VGND VPWR VPWR dadda_fa_5_10_1/A dadda_ha_4_9_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$1210 U$$525/A1 U$$1230/A2 U$$2171/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1211/A
+ sky130_fd_sc_hd__a22o_1
XU$$1221 U$$1221/A U$$1225/B VGND VGND VPWR VPWR U$$1221/X sky130_fd_sc_hd__xor2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1232 U$$1232/A VGND VGND VPWR VPWR U$$1232/Y sky130_fd_sc_hd__inv_1
XFILLER_44_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1243 U$$8/B1 U$$1279/A2 U$$12/A1 U$$1279/B2 VGND VGND VPWR VPWR U$$1244/A sky130_fd_sc_hd__a22o_1
XFILLER_50_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1254 U$$1254/A U$$1292/B VGND VGND VPWR VPWR U$$1254/X sky130_fd_sc_hd__xor2_1
XU$$1265 U$$854/A1 U$$1295/A2 U$$993/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1266/A sky130_fd_sc_hd__a22o_1
XFILLER_206_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1276 U$$1276/A U$$1280/B VGND VGND VPWR VPWR U$$1276/X sky130_fd_sc_hd__xor2_1
XU$$1287 U$$463/B1 U$$1323/A2 U$$330/A1 U$$1323/B2 VGND VGND VPWR VPWR U$$1288/A sky130_fd_sc_hd__a22o_1
XFILLER_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XU$$1298 U$$1298/A U$$1310/B VGND VGND VPWR VPWR U$$1298/X sky130_fd_sc_hd__xor2_1
XFILLER_175_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1028 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_84_1 dadda_fa_5_84_1/A dadda_fa_5_84_1/B dadda_fa_5_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_85_0/B dadda_fa_7_84_0/A sky130_fd_sc_hd__fa_2
XFILLER_117_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_77_0 dadda_fa_5_77_0/A dadda_fa_5_77_0/B dadda_fa_5_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_78_0/A dadda_fa_6_77_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_176_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_76_8 dadda_fa_1_76_8/A dadda_fa_1_76_8/B dadda_fa_1_76_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_77_3/A dadda_fa_3_76_0/A sky130_fd_sc_hd__fa_2
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_7 dadda_fa_1_69_7/A dadda_fa_1_69_7/B dadda_fa_1_69_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_2/CIN dadda_fa_2_69_5/CIN sky130_fd_sc_hd__fa_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3190 U$$3190/A U$$3236/B VGND VGND VPWR VPWR U$$3190/X sky130_fd_sc_hd__xor2_1
XFILLER_50_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_95_0 U$$2191/Y U$$2325/X U$$2458/X VGND VGND VPWR VPWR dadda_fa_2_96_5/CIN
+ dadda_fa_3_95_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_100_3 dadda_fa_3_100_3/A dadda_fa_3_100_3/B dadda_fa_3_100_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_1/B dadda_fa_4_100_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_2_108_0 dadda_ha_2_108_0/A U$$3149/X VGND VGND VPWR VPWR dadda_fa_4_109_0/A
+ dadda_fa_4_108_0/A sky130_fd_sc_hd__ha_1
XTAP_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$451 final_adder.U$$274/B final_adder.U$$658/B final_adder.U$$165/X
+ VGND VGND VPWR VPWR final_adder.U$$660/B sky130_fd_sc_hd__a21o_1
XTAP_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_622_ _623_/CLK _622_/D VGND VGND VPWR VPWR _622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$301 U$$301/A U$$309/B VGND VGND VPWR VPWR U$$301/X sky130_fd_sc_hd__xor2_1
XFILLER_18_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_107_0 dadda_fa_6_107_0/A dadda_fa_6_107_0/B dadda_fa_6_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_108_0/B dadda_fa_7_107_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$473 final_adder.U$$296/B final_adder.U$$702/B final_adder.U$$209/X
+ VGND VGND VPWR VPWR final_adder.U$$704/B sky130_fd_sc_hd__a21o_1
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$312 U$$449/A1 U$$318/A2 U$$449/B1 U$$318/B2 VGND VGND VPWR VPWR U$$313/A sky130_fd_sc_hd__a22o_1
XTAP_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$323 U$$323/A U$$335/B VGND VGND VPWR VPWR U$$323/X sky130_fd_sc_hd__xor2_1
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$495 final_adder.U$$252/X final_adder.U$$746/B final_adder.U$$253/X
+ VGND VGND VPWR VPWR final_adder.U$$748/B sky130_fd_sc_hd__a21o_2
XU$$334 U$$334/A1 U$$334/A2 U$$334/B1 U$$334/B2 VGND VGND VPWR VPWR U$$335/A sky130_fd_sc_hd__a22o_1
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$345 U$$345/A U$$351/B VGND VGND VPWR VPWR U$$345/X sky130_fd_sc_hd__xor2_1
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_553_ _558_/CLK _553_/D VGND VGND VPWR VPWR _553_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$356 U$$493/A1 U$$398/A2 U$$358/A1 U$$398/B2 VGND VGND VPWR VPWR U$$357/A sky130_fd_sc_hd__a22o_1
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_27_3 dadda_fa_3_27_3/A dadda_fa_3_27_3/B dadda_fa_3_27_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_28_1/B dadda_fa_4_27_2/CIN sky130_fd_sc_hd__fa_1
XU$$367 U$$367/A U$$410/A VGND VGND VPWR VPWR U$$367/X sky130_fd_sc_hd__xor2_1
XFILLER_199_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$378 U$$650/B1 U$$384/A2 U$$515/B1 U$$384/B2 VGND VGND VPWR VPWR U$$379/A sky130_fd_sc_hd__a22o_1
XFILLER_83_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$389 U$$389/A U$$393/B VGND VGND VPWR VPWR U$$389/X sky130_fd_sc_hd__xor2_1
X_484_ _484_/CLK _484_/D VGND VGND VPWR VPWR _484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_94_0 dadda_fa_6_94_0/A dadda_fa_6_94_0/B dadda_fa_6_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_95_0/B dadda_fa_7_94_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_185_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1201 U$$4105/A1 VGND VGND VPWR VPWR U$$406/A1 sky130_fd_sc_hd__buf_4
XFILLER_201_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1212 U$$2459/A1 VGND VGND VPWR VPWR U$$952/A1 sky130_fd_sc_hd__buf_6
Xrepeater1223 _612_/Q VGND VGND VPWR VPWR U$$3005/A1 sky130_fd_sc_hd__buf_6
XFILLER_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1234 U$$2314/B1 VGND VGND VPWR VPWR U$$946/A1 sky130_fd_sc_hd__buf_8
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1245 U$$3273/A1 VGND VGND VPWR VPWR U$$4506/A1 sky130_fd_sc_hd__buf_4
Xrepeater1256 U$$2858/A1 VGND VGND VPWR VPWR U$$253/B1 sky130_fd_sc_hd__buf_6
XFILLER_114_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1267 U$$4361/B1 VGND VGND VPWR VPWR U$$938/A1 sky130_fd_sc_hd__buf_4
Xrepeater1278 U$$4087/A1 VGND VGND VPWR VPWR U$$4498/A1 sky130_fd_sc_hd__buf_4
XFILLER_107_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1289 _604_/Q VGND VGND VPWR VPWR U$$3674/A1 sky130_fd_sc_hd__buf_4
XFILLER_141_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$890 U$$66/B1 U$$928/A2 U$$890/B1 U$$928/B2 VGND VGND VPWR VPWR U$$891/A sky130_fd_sc_hd__a22o_1
XU$$1040 U$$1040/A U$$1040/B VGND VGND VPWR VPWR U$$1040/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1051 U$$229/A1 U$$1093/A2 U$$368/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1052/A sky130_fd_sc_hd__a22o_1
XU$$1062 U$$1062/A U$$996/B VGND VGND VPWR VPWR U$$1062/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1073 U$$4224/A1 U$$963/X U$$527/A1 U$$964/X VGND VGND VPWR VPWR U$$1074/A sky130_fd_sc_hd__a22o_1
XU$$1084 U$$1084/A U$$1095/A VGND VGND VPWR VPWR U$$1084/X sky130_fd_sc_hd__xor2_1
XU$$1095 U$$1095/A VGND VGND VPWR VPWR U$$1095/Y sky130_fd_sc_hd__inv_1
XFILLER_149_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3157_1747 VGND VGND VPWR VPWR U$$3157_1747/HI U$$3157/A1 sky130_fd_sc_hd__conb_1
XFILLER_177_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_978 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_81_6 U$$3627/X U$$3760/X U$$3893/X VGND VGND VPWR VPWR dadda_fa_2_82_3/A
+ dadda_fa_2_81_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_171_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_74_5 U$$3746/X U$$3879/X U$$4012/X VGND VGND VPWR VPWR dadda_fa_2_75_2/A
+ dadda_fa_2_74_5/A sky130_fd_sc_hd__fa_1
XFILLER_98_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_4 U$$4131/X U$$4264/X U$$4397/X VGND VGND VPWR VPWR dadda_fa_2_68_1/CIN
+ dadda_fa_2_67_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_37_2 dadda_fa_4_37_2/A dadda_fa_4_37_2/B dadda_fa_4_37_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/CIN dadda_fa_5_37_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1020 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_842 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_63_5 U$$2128/X U$$2261/X VGND VGND VPWR VPWR dadda_fa_1_64_7/A dadda_fa_2_63_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_123_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_62_3 U$$1328/X U$$1461/X U$$1594/X VGND VGND VPWR VPWR dadda_fa_1_63_6/B
+ dadda_fa_1_62_8/B sky130_fd_sc_hd__fa_1
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3904 U$$4176/B1 U$$3968/A2 U$$4180/A1 U$$3968/B2 VGND VGND VPWR VPWR U$$3905/A
+ sky130_fd_sc_hd__a22o_1
XU$$3915 U$$3915/A U$$3917/B VGND VGND VPWR VPWR U$$3915/X sky130_fd_sc_hd__xor2_1
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3926 _593_/Q U$$3932/A2 U$$4337/B1 U$$3932/B2 VGND VGND VPWR VPWR U$$3927/A sky130_fd_sc_hd__a22o_1
XFILLER_64_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3937 U$$3937/A U$$3943/B VGND VGND VPWR VPWR U$$3937/X sky130_fd_sc_hd__xor2_1
XFILLER_206_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3948 U$$4494/B1 U$$3958/A2 U$$4498/A1 U$$3958/B2 VGND VGND VPWR VPWR U$$3949/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$270 final_adder.U$$270/A final_adder.U$$270/B VGND VGND VPWR VPWR
+ final_adder.U$$326/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$281 final_adder.U$$280/A final_adder.U$$177/X final_adder.U$$179/X
+ VGND VGND VPWR VPWR final_adder.U$$281/X sky130_fd_sc_hd__a21o_1
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_32_1 dadda_fa_3_32_1/A dadda_fa_3_32_1/B dadda_fa_3_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_0/CIN dadda_fa_4_32_2/A sky130_fd_sc_hd__fa_2
XU$$120 U$$942/A1 U$$128/A2 U$$942/B1 U$$128/B2 VGND VGND VPWR VPWR U$$121/A sky130_fd_sc_hd__a22o_1
X_605_ _613_/CLK _605_/D VGND VGND VPWR VPWR _605_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$292 final_adder.U$$292/A final_adder.U$$292/B VGND VGND VPWR VPWR
+ final_adder.U$$338/B sky130_fd_sc_hd__and2_1
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3959 U$$3959/A U$$3965/B VGND VGND VPWR VPWR U$$3959/X sky130_fd_sc_hd__xor2_1
XU$$131 U$$131/A U$$2/A VGND VGND VPWR VPWR U$$131/X sky130_fd_sc_hd__xor2_1
XFILLER_206_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$142 U$$140/B U$$2/A _618_/Q U$$137/Y VGND VGND VPWR VPWR U$$142/X sky130_fd_sc_hd__a22o_1
XFILLER_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$153 U$$16/A1 U$$181/A2 U$$18/A1 U$$181/B2 VGND VGND VPWR VPWR U$$154/A sky130_fd_sc_hd__a22o_1
XFILLER_18_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$164 U$$164/A U$$190/B VGND VGND VPWR VPWR U$$164/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_25_0 U$$722/X U$$855/X U$$988/X VGND VGND VPWR VPWR dadda_fa_4_26_0/B
+ dadda_fa_4_25_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_60_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$175 U$$997/A1 U$$175/A2 U$$40/A1 U$$175/B2 VGND VGND VPWR VPWR U$$176/A sky130_fd_sc_hd__a22o_1
X_536_ _538_/CLK _536_/D VGND VGND VPWR VPWR _536_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$186 U$$186/A U$$232/B VGND VGND VPWR VPWR U$$186/X sky130_fd_sc_hd__xor2_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$197 U$$60/A1 U$$263/A2 U$$62/A1 U$$263/B2 VGND VGND VPWR VPWR U$$198/A sky130_fd_sc_hd__a22o_1
XFILLER_207_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_467_ _467_/CLK _467_/D VGND VGND VPWR VPWR _467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_398_ _615_/CLK _398_/D VGND VGND VPWR VPWR _398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_91_5 dadda_fa_2_91_5/A dadda_fa_2_91_5/B dadda_fa_2_91_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_92_2/A dadda_fa_4_91_0/A sky130_fd_sc_hd__fa_1
XFILLER_12_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1020 _655_/Q VGND VGND VPWR VPWR U$$2739/A sky130_fd_sc_hd__buf_6
XFILLER_127_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1031 U$$2466/A VGND VGND VPWR VPWR U$$2465/A sky130_fd_sc_hd__buf_6
XFILLER_127_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1042 U$$2309/B VGND VGND VPWR VPWR U$$2303/B sky130_fd_sc_hd__buf_8
XFILLER_86_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1053 U$$2186/B VGND VGND VPWR VPWR U$$2191/A sky130_fd_sc_hd__buf_6
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2061_1729 VGND VGND VPWR VPWR U$$2061_1729/HI U$$2061/A1 sky130_fd_sc_hd__conb_1
Xrepeater1064 _645_/Q VGND VGND VPWR VPWR U$$2003/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_84_4 dadda_fa_2_84_4/A dadda_fa_2_84_4/B dadda_fa_2_84_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/CIN dadda_fa_3_84_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1075 _641_/Q VGND VGND VPWR VPWR U$$1737/B sky130_fd_sc_hd__buf_6
XFILLER_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1086 _639_/Q VGND VGND VPWR VPWR U$$1642/B sky130_fd_sc_hd__buf_6
Xrepeater1097 U$$1501/B VGND VGND VPWR VPWR U$$1487/B sky130_fd_sc_hd__buf_6
XFILLER_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_77_3 dadda_fa_2_77_3/A dadda_fa_2_77_3/B dadda_fa_2_77_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/B dadda_fa_3_77_3/B sky130_fd_sc_hd__fa_1
XFILLER_68_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_47_1 dadda_fa_5_47_1/A dadda_fa_5_47_1/B dadda_fa_5_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_48_0/B dadda_fa_7_47_0/A sky130_fd_sc_hd__fa_1
XFILLER_96_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_100_2 U$$3266/X U$$3399/X U$$3532/X VGND VGND VPWR VPWR dadda_fa_3_101_2/A
+ dadda_fa_3_100_3/B sky130_fd_sc_hd__fa_1
XFILLER_24_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_121_1 dadda_fa_5_121_1/A dadda_fa_5_121_1/B dadda_fa_5_121_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_122_0/B dadda_fa_7_121_0/A sky130_fd_sc_hd__fa_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_114_0 dadda_fa_5_114_0/A dadda_fa_5_114_0/B dadda_fa_5_114_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_115_0/A dadda_fa_6_114_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_165_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_2_0_clk/X sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_1_72_2 U$$2811/X U$$2944/X U$$3077/X VGND VGND VPWR VPWR dadda_fa_2_73_1/A
+ dadda_fa_2_72_4/A sky130_fd_sc_hd__fa_1
XFILLER_58_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_65_1 U$$2930/X U$$3063/X U$$3196/X VGND VGND VPWR VPWR dadda_fa_2_66_0/CIN
+ dadda_fa_2_65_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_42_0 dadda_fa_4_42_0/A dadda_fa_4_42_0/B dadda_fa_4_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/A dadda_fa_5_42_1/A sky130_fd_sc_hd__fa_1
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_58_0 U$$1586/X U$$1719/X U$$1852/X VGND VGND VPWR VPWR dadda_fa_2_59_0/B
+ dadda_fa_2_58_3/B sky130_fd_sc_hd__fa_1
XFILLER_101_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1809 U$$848/B1 U$$1851/A2 U$$715/A1 U$$1851/B2 VGND VGND VPWR VPWR U$$1810/A sky130_fd_sc_hd__a22o_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_321_ _451_/CLK _321_/D VGND VGND VPWR VPWR _321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_52 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_252_ _253_/CLK _252_/D VGND VGND VPWR VPWR _252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_183_ _189_/CLK _183_/D VGND VGND VPWR VPWR _183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_446 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_94_3 dadda_fa_3_94_3/A dadda_fa_3_94_3/B dadda_fa_3_94_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_1/B dadda_fa_4_94_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_129_83 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_87_2 dadda_fa_3_87_2/A dadda_fa_3_87_2/B dadda_fa_3_87_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_1/A dadda_fa_4_87_2/B sky130_fd_sc_hd__fa_1
XFILLER_151_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_54_1 U$$514/X U$$647/X VGND VGND VPWR VPWR dadda_fa_1_55_8/B dadda_fa_2_54_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_57_0 dadda_fa_6_57_0/A dadda_fa_6_57_0/B dadda_fa_6_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_58_0/B dadda_fa_7_57_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_81_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater709 U$$3841/X VGND VGND VPWR VPWR U$$3968/B2 sky130_fd_sc_hd__buf_6
XU$$4402 U$$4402/A1 U$$4388/X U$$4402/B1 U$$4438/B2 VGND VGND VPWR VPWR U$$4403/A
+ sky130_fd_sc_hd__a22o_1
XU$$4413 U$$4413/A U$$4413/B VGND VGND VPWR VPWR U$$4413/X sky130_fd_sc_hd__xor2_1
XU$$4424 _568_/Q U$$4388/X U$$4426/A1 U$$4454/B2 VGND VGND VPWR VPWR U$$4425/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_0_60_0 U$$127/X U$$260/X U$$393/X VGND VGND VPWR VPWR dadda_fa_1_61_6/A
+ dadda_fa_1_60_7/CIN sky130_fd_sc_hd__fa_1
XU$$4435 U$$4435/A U$$4435/B VGND VGND VPWR VPWR U$$4435/X sky130_fd_sc_hd__xor2_1
XU$$4446 _579_/Q U$$4388/X U$$4446/B1 U$$4468/B2 VGND VGND VPWR VPWR U$$4447/A sky130_fd_sc_hd__a22o_1
XFILLER_77_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3701 U$$3835/A VGND VGND VPWR VPWR U$$3701/Y sky130_fd_sc_hd__inv_1
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3712 U$$3712/A U$$3764/B VGND VGND VPWR VPWR U$$3712/X sky130_fd_sc_hd__xor2_1
XU$$4457 U$$4457/A U$$4457/B VGND VGND VPWR VPWR U$$4457/X sky130_fd_sc_hd__xor2_1
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_116_2 input147/X dadda_fa_4_116_2/B dadda_ha_3_116_0/SUM VGND VGND VPWR
+ VPWR dadda_fa_5_117_0/CIN dadda_fa_5_116_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3723 _560_/Q U$$3833/A2 U$$4136/A1 U$$3833/B2 VGND VGND VPWR VPWR U$$3724/A sky130_fd_sc_hd__a22o_1
XU$$4468 U$$4468/A1 U$$4388/X U$$4470/A1 U$$4468/B2 VGND VGND VPWR VPWR U$$4469/A
+ sky130_fd_sc_hd__a22o_1
XU$$3734 U$$3734/A U$$3816/B VGND VGND VPWR VPWR U$$3734/X sky130_fd_sc_hd__xor2_1
XU$$4479 U$$4479/A U$$4479/B VGND VGND VPWR VPWR U$$4479/X sky130_fd_sc_hd__xor2_1
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3745 U$$4154/B1 U$$3785/A2 U$$4156/B1 U$$3785/B2 VGND VGND VPWR VPWR U$$3746/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3756 U$$3756/A U$$3760/B VGND VGND VPWR VPWR U$$3756/X sky130_fd_sc_hd__xor2_1
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_109_1 dadda_fa_4_109_1/A dadda_fa_4_109_1/B dadda_fa_4_109_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/B dadda_fa_5_109_1/B sky130_fd_sc_hd__fa_1
XU$$3767 U$$3902/B1 U$$3823/A2 U$$3769/A1 U$$3823/B2 VGND VGND VPWR VPWR U$$3768/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3778 U$$3778/A _671_/Q VGND VGND VPWR VPWR U$$3778/X sky130_fd_sc_hd__xor2_1
XU$$3789 _593_/Q U$$3795/A2 U$$3789/B1 U$$3795/B2 VGND VGND VPWR VPWR U$$3790/A sky130_fd_sc_hd__a22o_1
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_360 U$$2981/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_371 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_519_ _519_/CLK _519_/D VGND VGND VPWR VPWR _519_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_382 _640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_393 U$$1478/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_82_1 dadda_fa_2_82_1/A dadda_fa_2_82_1/B dadda_fa_2_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_0/CIN dadda_fa_3_82_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_75_0 dadda_fa_2_75_0/A dadda_fa_2_75_0/B dadda_fa_2_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_0/B dadda_fa_3_75_2/B sky130_fd_sc_hd__fa_1
XFILLER_130_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_51_7 U$$2902/X U$$3035/X U$$3168/X VGND VGND VPWR VPWR dadda_fa_2_52_2/CIN
+ dadda_fa_2_51_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_84_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1025 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_97_1 dadda_fa_4_97_1/A dadda_fa_4_97_1/B dadda_fa_4_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/B dadda_fa_5_97_1/B sky130_fd_sc_hd__fa_1
XFILLER_30_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_74_0 dadda_fa_7_74_0/A dadda_fa_7_74_0/B dadda_fa_7_74_0/CIN VGND VGND
+ VPWR VPWR _499_/D _370_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_2_104_0_1864 VGND VGND VPWR VPWR dadda_fa_2_104_0/A dadda_fa_2_104_0_1864/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_124_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_23 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3008 U$$3008/A U$$3008/B VGND VGND VPWR VPWR U$$3008/X sky130_fd_sc_hd__xor2_1
XU$$3019 U$$3017/B U$$3014/A _660_/Q U$$3014/Y VGND VGND VPWR VPWR U$$3019/X sky130_fd_sc_hd__a22o_1
XU$$2307 U$$2307/A U$$2309/B VGND VGND VPWR VPWR U$$2307/X sky130_fd_sc_hd__xor2_1
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2318 _611_/Q U$$2318/A2 U$$2318/B1 U$$2318/B2 VGND VGND VPWR VPWR U$$2319/A sky130_fd_sc_hd__a22o_1
XU$$2329 _649_/Q VGND VGND VPWR VPWR U$$2329/Y sky130_fd_sc_hd__inv_1
XU$$1606 U$$1606/A U$$1642/B VGND VGND VPWR VPWR U$$1606/X sky130_fd_sc_hd__xor2_1
XU$$1617 U$$382/B1 U$$1627/A2 U$$384/B1 U$$1627/B2 VGND VGND VPWR VPWR U$$1618/A sky130_fd_sc_hd__a22o_1
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1628 U$$1628/A U$$1628/B VGND VGND VPWR VPWR U$$1628/X sky130_fd_sc_hd__xor2_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1639 U$$678/B1 U$$1511/X U$$545/A1 U$$1512/X VGND VGND VPWR VPWR U$$1640/A sky130_fd_sc_hd__a22o_1
XFILLER_203_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_304_ _442_/CLK _304_/D VGND VGND VPWR VPWR _304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_235_ _503_/CLK _235_/D VGND VGND VPWR VPWR _235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_92_0 dadda_fa_3_92_0/A dadda_fa_3_92_0/B dadda_fa_3_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_0/B dadda_fa_4_92_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_155_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater506 U$$3148/A2 VGND VGND VPWR VPWR U$$3110/A2 sky130_fd_sc_hd__buf_8
XFILLER_78_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater517 U$$2881/X VGND VGND VPWR VPWR U$$3005/A2 sky130_fd_sc_hd__buf_4
XU$$4210 U$$4484/A1 U$$4244/A2 U$$4486/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4211/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater528 U$$2832/A2 VGND VGND VPWR VPWR U$$2812/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_54_5 dadda_fa_2_54_5/A dadda_fa_2_54_5/B dadda_fa_2_54_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_2/A dadda_fa_4_54_0/A sky130_fd_sc_hd__fa_1
Xrepeater539 U$$2729/A2 VGND VGND VPWR VPWR U$$2687/A2 sky130_fd_sc_hd__buf_4
XFILLER_133_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4221 U$$4221/A U$$4246/A VGND VGND VPWR VPWR U$$4221/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_121_0 U$$3972/Y U$$4106/X U$$4239/X VGND VGND VPWR VPWR dadda_fa_5_122_1/B
+ dadda_fa_5_121_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4232 U$$4369/A1 U$$4238/A2 U$$4369/B1 U$$4238/B2 VGND VGND VPWR VPWR U$$4233/A
+ sky130_fd_sc_hd__a22o_1
XU$$4243 U$$4243/A U$$4246/A VGND VGND VPWR VPWR U$$4243/X sky130_fd_sc_hd__xor2_1
XFILLER_92_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4254 U$$4254/A U$$4298/B VGND VGND VPWR VPWR U$$4254/X sky130_fd_sc_hd__xor2_1
XU$$3520 U$$3520/A U$$3520/B VGND VGND VPWR VPWR U$$3520/X sky130_fd_sc_hd__xor2_1
XU$$4265 U$$4402/A1 U$$4347/A2 _558_/Q U$$4347/B2 VGND VGND VPWR VPWR U$$4266/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_47_4 dadda_fa_2_47_4/A dadda_fa_2_47_4/B dadda_fa_2_47_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/CIN dadda_fa_3_47_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_207_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3531 U$$3805/A1 U$$3531/A2 U$$3805/B1 U$$3531/B2 VGND VGND VPWR VPWR U$$3532/A
+ sky130_fd_sc_hd__a22o_1
XU$$4276 U$$4276/A U$$4296/B VGND VGND VPWR VPWR U$$4276/X sky130_fd_sc_hd__xor2_1
XFILLER_77_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3542 U$$3542/A _667_/Q VGND VGND VPWR VPWR U$$3542/X sky130_fd_sc_hd__xor2_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4287 U$$4287/A1 U$$4311/A2 U$$4426/A1 U$$4311/B2 VGND VGND VPWR VPWR U$$4288/A
+ sky130_fd_sc_hd__a22o_1
XU$$3553 U$$4512/A1 U$$3555/A2 U$$4514/A1 U$$3555/B2 VGND VGND VPWR VPWR U$$3554/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4298 U$$4298/A U$$4298/B VGND VGND VPWR VPWR U$$4298/X sky130_fd_sc_hd__xor2_1
XU$$3564 _669_/Q VGND VGND VPWR VPWR U$$3564/Y sky130_fd_sc_hd__inv_1
XU$$3575 U$$3575/A U$$3613/B VGND VGND VPWR VPWR U$$3575/X sky130_fd_sc_hd__xor2_1
XFILLER_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2830 U$$2830/A1 U$$2832/A2 U$$229/A1 U$$2832/B2 VGND VGND VPWR VPWR U$$2831/A
+ sky130_fd_sc_hd__a22o_1
XU$$3586 U$$4408/A1 U$$3628/A2 U$$4136/A1 U$$3628/B2 VGND VGND VPWR VPWR U$$3587/A
+ sky130_fd_sc_hd__a22o_1
XU$$2841 U$$2841/A U$$2843/B VGND VGND VPWR VPWR U$$2841/X sky130_fd_sc_hd__xor2_1
XFILLER_80_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2852 U$$3124/B1 U$$2856/A2 U$$2991/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2853/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_448 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3597 U$$3597/A U$$3637/B VGND VGND VPWR VPWR U$$3597/X sky130_fd_sc_hd__xor2_1
XFILLER_206_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2863 U$$2863/A _657_/Q VGND VGND VPWR VPWR U$$2863/X sky130_fd_sc_hd__xor2_1
XU$$2874 U$$3285/A1 U$$2874/A2 U$$2874/B1 U$$2874/B2 VGND VGND VPWR VPWR U$$2875/A
+ sky130_fd_sc_hd__a22o_1
XU$$2885 U$$3157/B1 U$$2929/A2 U$$3022/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2886/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2896 U$$2896/A U$$2944/B VGND VGND VPWR VPWR U$$2896/X sky130_fd_sc_hd__xor2_1
XFILLER_205_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_190 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_984 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$708 U$$708/A U$$726/B VGND VGND VPWR VPWR U$$708/X sky130_fd_sc_hd__xor2_1
XFILLER_56_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$719 U$$993/A1 U$$759/A2 U$$719/B1 U$$759/B2 VGND VGND VPWR VPWR U$$720/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_42_3 U$$1288/X U$$1421/X U$$1554/X VGND VGND VPWR VPWR dadda_fa_2_43_4/A
+ dadda_fa_2_42_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_12_1 U$$430/X U$$563/X U$$696/X VGND VGND VPWR VPWR dadda_fa_5_13_0/B
+ dadda_fa_5_12_1/B sky130_fd_sc_hd__fa_1
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1608 U$$3181/B1 VGND VGND VPWR VPWR U$$4140/B1 sky130_fd_sc_hd__buf_8
XFILLER_137_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1619 _563_/Q VGND VGND VPWR VPWR U$$4140/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_109_0 U$$3150/Y U$$3284/X U$$3417/X VGND VGND VPWR VPWR dadda_fa_4_110_0/B
+ dadda_fa_4_109_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_57_3 dadda_fa_3_57_3/A dadda_fa_3_57_3/B dadda_fa_3_57_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_1/B dadda_fa_4_57_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2104 U$$2104/A U$$2110/B VGND VGND VPWR VPWR U$$2104/X sky130_fd_sc_hd__xor2_1
XFILLER_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_724 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2115 U$$4031/B1 U$$2115/A2 U$$3213/A1 U$$2115/B2 VGND VGND VPWR VPWR U$$2116/A
+ sky130_fd_sc_hd__a22o_1
XU$$2126 U$$2126/A U$$2136/B VGND VGND VPWR VPWR U$$2126/X sky130_fd_sc_hd__xor2_1
XU$$2137 U$$3505/B1 U$$2059/X U$$3372/A1 U$$2060/X VGND VGND VPWR VPWR U$$2138/A sky130_fd_sc_hd__a22o_1
XU$$1403 U$$1403/A U$$1443/B VGND VGND VPWR VPWR U$$1403/X sky130_fd_sc_hd__xor2_1
XU$$2148 U$$2148/A U$$2170/B VGND VGND VPWR VPWR U$$2148/X sky130_fd_sc_hd__xor2_1
XFILLER_188_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2159 U$$2431/B1 U$$2189/A2 U$$3255/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2160/A
+ sky130_fd_sc_hd__a22o_1
XU$$1414 U$$866/A1 U$$1428/A2 U$$866/B1 U$$1428/B2 VGND VGND VPWR VPWR U$$1415/A sky130_fd_sc_hd__a22o_1
XU$$1425 U$$1425/A U$$1425/B VGND VGND VPWR VPWR U$$1425/X sky130_fd_sc_hd__xor2_1
XFILLER_76_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1436 U$$614/A1 U$$1442/A2 U$$614/B1 U$$1442/B2 VGND VGND VPWR VPWR U$$1437/A sky130_fd_sc_hd__a22o_1
XFILLER_16_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1447 U$$1447/A U$$1487/B VGND VGND VPWR VPWR U$$1447/X sky130_fd_sc_hd__xor2_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1458 U$$88/A1 U$$1458/A2 U$$90/A1 U$$1458/B2 VGND VGND VPWR VPWR U$$1459/A sky130_fd_sc_hd__a22o_1
XU$$3294_1749 VGND VGND VPWR VPWR U$$3294_1749/HI U$$3294/A1 sky130_fd_sc_hd__conb_1
XU$$1469 U$$1469/A U$$1475/B VGND VGND VPWR VPWR U$$1469/X sky130_fd_sc_hd__xor2_1
XFILLER_35_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_218_ _351_/CLK _218_/D VGND VGND VPWR VPWR _218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_52_2 dadda_fa_2_52_2/A dadda_fa_2_52_2/B dadda_fa_2_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/A dadda_fa_3_52_3/A sky130_fd_sc_hd__fa_1
XFILLER_38_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4040 U$$4040/A U$$4072/B VGND VGND VPWR VPWR U$$4040/X sky130_fd_sc_hd__xor2_1
XFILLER_38_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4051 U$$4051/A1 U$$4061/A2 U$$4053/A1 U$$4061/B2 VGND VGND VPWR VPWR U$$4052/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_45_1 U$$2757/X U$$2890/X U$$3023/X VGND VGND VPWR VPWR dadda_fa_3_46_0/CIN
+ dadda_fa_3_45_2/CIN sky130_fd_sc_hd__fa_1
XU$$4062 U$$4062/A U$$4070/B VGND VGND VPWR VPWR U$$4062/X sky130_fd_sc_hd__xor2_1
XFILLER_38_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4073 U$$4208/B1 U$$3977/X U$$4486/A1 U$$3978/X VGND VGND VPWR VPWR U$$4074/A sky130_fd_sc_hd__a22o_1
XU$$4084 U$$4084/A U$$4084/B VGND VGND VPWR VPWR U$$4084/X sky130_fd_sc_hd__xor2_1
XFILLER_81_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3350 U$$3624/A1 U$$3404/A2 U$$3352/A1 U$$3404/B2 VGND VGND VPWR VPWR U$$3351/A
+ sky130_fd_sc_hd__a22o_1
XU$$4095 U$$805/B1 U$$4095/A2 U$$4369/B1 U$$4105/B2 VGND VGND VPWR VPWR U$$4096/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_22_0 dadda_fa_5_22_0/A dadda_fa_5_22_0/B dadda_fa_5_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_23_0/A dadda_fa_6_22_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_38_0 U$$1147/X U$$1280/X U$$1413/X VGND VGND VPWR VPWR dadda_fa_3_39_0/B
+ dadda_fa_3_38_2/B sky130_fd_sc_hd__fa_1
XU$$3361 U$$3361/A U$$3363/B VGND VGND VPWR VPWR U$$3361/X sky130_fd_sc_hd__xor2_1
XFILLER_19_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3372 U$$3372/A1 U$$3418/A2 U$$3374/A1 U$$3418/B2 VGND VGND VPWR VPWR U$$3373/A
+ sky130_fd_sc_hd__a22o_1
XU$$3383 U$$3383/A U$$3397/B VGND VGND VPWR VPWR U$$3383/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3394 _601_/Q U$$3402/A2 _602_/Q U$$3402/B2 VGND VGND VPWR VPWR U$$3395/A sky130_fd_sc_hd__a22o_1
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2660 U$$2660/A U$$2664/B VGND VGND VPWR VPWR U$$2660/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2671 U$$3902/B1 U$$2707/A2 U$$3769/A1 U$$2707/B2 VGND VGND VPWR VPWR U$$2672/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2682 U$$2682/A U$$2698/B VGND VGND VPWR VPWR U$$2682/X sky130_fd_sc_hd__xor2_1
XU$$2693 U$$2830/A1 U$$2733/A2 U$$3789/B1 U$$2733/B2 VGND VGND VPWR VPWR U$$2694/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1970 U$$3751/A1 U$$1976/A2 U$$3753/A1 U$$1976/B2 VGND VGND VPWR VPWR U$$1971/A
+ sky130_fd_sc_hd__a22o_1
XU$$1981 U$$1981/A U$$2029/B VGND VGND VPWR VPWR U$$1981/X sky130_fd_sc_hd__xor2_1
XFILLER_179_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1992 U$$759/A1 U$$1922/X U$$624/A1 U$$1923/X VGND VGND VPWR VPWR U$$1993/A sky130_fd_sc_hd__a22o_1
XFILLER_178_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_67_2 dadda_fa_4_67_2/A dadda_fa_4_67_2/B dadda_fa_4_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/CIN dadda_fa_5_67_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput106 b[47] VGND VGND VPWR VPWR _599_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput117 b[57] VGND VGND VPWR VPWR _609_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput128 b[9] VGND VGND VPWR VPWR _561_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput139 c[109] VGND VGND VPWR VPWR input139/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_37_0 dadda_fa_7_37_0/A dadda_fa_7_37_0/B dadda_fa_7_37_0/CIN VGND VGND
+ VPWR VPWR _462_/D _333_/D sky130_fd_sc_hd__fa_1
XTAP_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$611 final_adder.U$$738/A final_adder.U$$738/B final_adder.U$$611/B1
+ VGND VGND VPWR VPWR final_adder.U$$739/B sky130_fd_sc_hd__a21o_1
XFILLER_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$622 final_adder.U$$622/A final_adder.U$$622/B VGND VGND VPWR VPWR
+ _168_/D sky130_fd_sc_hd__xor2_1
XTAP_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$633 final_adder.U$$633/A final_adder.U$$633/B VGND VGND VPWR VPWR
+ _179_/D sky130_fd_sc_hd__xor2_4
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$644 final_adder.U$$644/A final_adder.U$$644/B VGND VGND VPWR VPWR
+ _190_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$655 final_adder.U$$655/A final_adder.U$$655/B VGND VGND VPWR VPWR
+ _201_/D sky130_fd_sc_hd__xor2_1
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$505 U$$914/B1 U$$517/A2 U$$916/B1 U$$517/B2 VGND VGND VPWR VPWR U$$506/A sky130_fd_sc_hd__a22o_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater870 U$$1375/X VGND VGND VPWR VPWR U$$1478/B2 sky130_fd_sc_hd__clkbuf_8
Xfinal_adder.U$$666 final_adder.U$$666/A final_adder.U$$666/B VGND VGND VPWR VPWR
+ _212_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$677 final_adder.U$$677/A final_adder.U$$677/B VGND VGND VPWR VPWR
+ _223_/D sky130_fd_sc_hd__xor2_1
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$516 U$$516/A U$$518/B VGND VGND VPWR VPWR U$$516/X sky130_fd_sc_hd__xor2_1
XFILLER_5_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_40_0 U$$87/X U$$220/X U$$353/X VGND VGND VPWR VPWR dadda_fa_2_41_3/CIN
+ dadda_fa_2_40_5/A sky130_fd_sc_hd__fa_1
Xrepeater881 U$$1176/B2 VGND VGND VPWR VPWR U$$1146/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$527 U$$527/A1 U$$415/X U$$938/B1 U$$416/X VGND VGND VPWR VPWR U$$528/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$688 final_adder.U$$688/A final_adder.U$$688/B VGND VGND VPWR VPWR
+ _234_/D sky130_fd_sc_hd__xor2_4
XFILLER_84_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater892 U$$98/B2 VGND VGND VPWR VPWR U$$84/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$699 final_adder.U$$699/A final_adder.U$$699/B VGND VGND VPWR VPWR
+ _245_/D sky130_fd_sc_hd__xor2_1
XU$$538 U$$538/A _623_/Q VGND VGND VPWR VPWR U$$538/X sky130_fd_sc_hd__xor2_1
XFILLER_99_1097 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_1056 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$549 _624_/Q VGND VGND VPWR VPWR U$$551/B sky130_fd_sc_hd__inv_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_90 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1095 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1405 U$$3096/A1 VGND VGND VPWR VPWR U$$82/A1 sky130_fd_sc_hd__buf_4
XFILLER_153_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1416 U$$4464/A1 VGND VGND VPWR VPWR U$$3642/A1 sky130_fd_sc_hd__buf_6
XFILLER_125_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1427 U$$76/A1 VGND VGND VPWR VPWR U$$898/A1 sky130_fd_sc_hd__buf_6
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1438 U$$4184/A1 VGND VGND VPWR VPWR U$$3362/A1 sky130_fd_sc_hd__buf_6
XFILLER_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1449 U$$4045/A1 VGND VGND VPWR VPWR U$$3769/B1 sky130_fd_sc_hd__buf_4
XFILLER_193_1038 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_62_1 dadda_fa_3_62_1/A dadda_fa_3_62_1/B dadda_fa_3_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_0/CIN dadda_fa_4_62_2/A sky130_fd_sc_hd__fa_1
XFILLER_97_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_55_0 dadda_fa_3_55_0/A dadda_fa_3_55_0/B dadda_fa_3_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_0/B dadda_fa_4_55_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1200 U$$926/A1 U$$1208/A2 U$$928/A1 U$$1208/B2 VGND VGND VPWR VPWR U$$1201/A sky130_fd_sc_hd__a22o_1
XU$$1211 U$$1211/A U$$1232/A VGND VGND VPWR VPWR U$$1211/X sky130_fd_sc_hd__xor2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1222 U$$948/A1 U$$1224/A2 U$$948/B1 U$$1224/B2 VGND VGND VPWR VPWR U$$1223/A sky130_fd_sc_hd__a22o_1
XU$$1233 _633_/Q VGND VGND VPWR VPWR U$$1233/Y sky130_fd_sc_hd__inv_1
XFILLER_204_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1244 U$$1244/A U$$1280/B VGND VGND VPWR VPWR U$$1244/X sky130_fd_sc_hd__xor2_1
XFILLER_44_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1255 U$$568/B1 U$$1291/A2 U$$435/A1 U$$1291/B2 VGND VGND VPWR VPWR U$$1256/A sky130_fd_sc_hd__a22o_1
XU$$1266 U$$1266/A U$$1296/B VGND VGND VPWR VPWR U$$1266/X sky130_fd_sc_hd__xor2_1
XFILLER_189_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1277 U$$44/A1 U$$1279/A2 U$$46/A1 U$$1279/B2 VGND VGND VPWR VPWR U$$1278/A sky130_fd_sc_hd__a22o_1
XU$$1288 U$$1288/A U$$1288/B VGND VGND VPWR VPWR U$$1288/X sky130_fd_sc_hd__xor2_1
XU$$1299 U$$749/B1 U$$1309/A2 U$$68/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1300/A sky130_fd_sc_hd__a22o_1
XFILLER_175_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_112_0 dadda_fa_7_112_0/A dadda_fa_7_112_0/B dadda_fa_7_112_0/CIN VGND
+ VGND VPWR VPWR _537_/D _408_/D sky130_fd_sc_hd__fa_1
XFILLER_102_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_77_1 dadda_fa_5_77_1/A dadda_fa_5_77_1/B dadda_fa_5_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_78_0/B dadda_fa_7_77_0/A sky130_fd_sc_hd__fa_1
XFILLER_144_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_8 dadda_fa_1_69_8/A dadda_fa_1_69_8/B dadda_fa_1_69_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_3/A dadda_fa_3_69_0/A sky130_fd_sc_hd__fa_2
XFILLER_26_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_359 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3180 U$$3180/A U$$3232/B VGND VGND VPWR VPWR U$$3180/X sky130_fd_sc_hd__xor2_1
XU$$3191 U$$3602/A1 U$$3235/A2 U$$3193/A1 U$$3235/B2 VGND VGND VPWR VPWR U$$3192/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_9_0 dadda_fa_6_9_0/A dadda_fa_6_9_0/B dadda_fa_6_9_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_10_0/B dadda_fa_7_9_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2490 U$$3584/B1 U$$2530/A2 U$$435/B1 U$$2530/B2 VGND VGND VPWR VPWR U$$2491/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4453_1805 VGND VGND VPWR VPWR U$$4453_1805/HI U$$4453/B sky130_fd_sc_hd__conb_1
XFILLER_190_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_72_0 dadda_fa_4_72_0/A dadda_fa_4_72_0/B dadda_fa_4_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/A dadda_fa_5_72_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_88_0 dadda_fa_1_88_0/A U$$1779/X U$$1912/X VGND VGND VPWR VPWR dadda_fa_2_89_3/B
+ dadda_fa_2_88_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$441 final_adder.U$$264/B final_adder.U$$638/B final_adder.U$$145/X
+ VGND VGND VPWR VPWR final_adder.U$$640/B sky130_fd_sc_hd__a21o_1
XTAP_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_621_ _624_/CLK _621_/D VGND VGND VPWR VPWR _621_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$463 final_adder.U$$286/B final_adder.U$$682/B final_adder.U$$189/X
+ VGND VGND VPWR VPWR final_adder.U$$684/B sky130_fd_sc_hd__a21o_1
XTAP_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$302 U$$302/A1 U$$334/A2 U$$989/A1 U$$334/B2 VGND VGND VPWR VPWR U$$303/A sky130_fd_sc_hd__a22o_1
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_584 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$313 U$$313/A U$$319/B VGND VGND VPWR VPWR U$$313/X sky130_fd_sc_hd__xor2_1
XFILLER_205_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$485 final_adder.U$$308/B final_adder.U$$726/B final_adder.U$$233/X
+ VGND VGND VPWR VPWR final_adder.U$$728/B sky130_fd_sc_hd__a21o_1
XU$$324 U$$733/B1 U$$334/A2 U$$600/A1 U$$334/B2 VGND VGND VPWR VPWR U$$325/A sky130_fd_sc_hd__a22o_1
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$335 U$$335/A U$$335/B VGND VGND VPWR VPWR U$$335/X sky130_fd_sc_hd__xor2_1
XFILLER_83_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_552_ _552_/CLK _552_/D VGND VGND VPWR VPWR _552_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$346 U$$72/A1 U$$350/A2 U$$74/A1 U$$350/B2 VGND VGND VPWR VPWR U$$347/A sky130_fd_sc_hd__a22o_1
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$357 U$$357/A U$$397/B VGND VGND VPWR VPWR U$$357/X sky130_fd_sc_hd__xor2_1
XFILLER_205_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$368 U$$368/A1 U$$392/A2 U$$96/A1 U$$392/B2 VGND VGND VPWR VPWR U$$369/A sky130_fd_sc_hd__a22o_1
XU$$379 U$$379/A U$$383/B VGND VGND VPWR VPWR U$$379/X sky130_fd_sc_hd__xor2_1
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_483_ _484_/CLK _483_/D VGND VGND VPWR VPWR _483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_87_0 dadda_fa_6_87_0/A dadda_fa_6_87_0/B dadda_fa_6_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_88_0/B dadda_fa_7_87_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1202 U$$678/B1 VGND VGND VPWR VPWR U$$4105/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1213 U$$3281/A1 VGND VGND VPWR VPWR U$$4514/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_201_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1224 _611_/Q VGND VGND VPWR VPWR U$$948/A1 sky130_fd_sc_hd__buf_6
XFILLER_154_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1235 U$$2999/B1 VGND VGND VPWR VPWR U$$2314/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1246 _609_/Q VGND VGND VPWR VPWR U$$3273/A1 sky130_fd_sc_hd__buf_6
XFILLER_181_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1257 U$$3132/A1 VGND VGND VPWR VPWR U$$392/A1 sky130_fd_sc_hd__buf_6
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1268 U$$4087/B1 VGND VGND VPWR VPWR U$$4361/B1 sky130_fd_sc_hd__buf_8
Xrepeater1279 U$$3539/A1 VGND VGND VPWR VPWR U$$4087/A1 sky130_fd_sc_hd__buf_4
XU$$1924_1727 VGND VGND VPWR VPWR U$$1924_1727/HI U$$1924/A1 sky130_fd_sc_hd__conb_1
XFILLER_80_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$880 U$$880/A1 U$$896/A2 U$$882/A1 U$$896/B2 VGND VGND VPWR VPWR U$$881/A sky130_fd_sc_hd__a22o_1
XFILLER_23_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1030 U$$1030/A U$$982/B VGND VGND VPWR VPWR U$$1030/X sky130_fd_sc_hd__xor2_1
XU$$891 U$$891/A U$$935/B VGND VGND VPWR VPWR U$$891/X sky130_fd_sc_hd__xor2_1
XFILLER_50_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1041 U$$80/B1 U$$1089/A2 U$$906/A1 U$$1089/B2 VGND VGND VPWR VPWR U$$1042/A sky130_fd_sc_hd__a22o_1
XFILLER_189_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1052 U$$1052/A U$$1095/A VGND VGND VPWR VPWR U$$1052/X sky130_fd_sc_hd__xor2_1
XFILLER_189_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1063 U$$926/A1 U$$1065/A2 U$$928/A1 U$$1065/B2 VGND VGND VPWR VPWR U$$1064/A sky130_fd_sc_hd__a22o_1
XFILLER_91_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1074 U$$1074/A U$$1078/B VGND VGND VPWR VPWR U$$1074/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1085 U$$948/A1 U$$1093/A2 U$$948/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1086/A sky130_fd_sc_hd__a22o_1
XU$$1096 _631_/Q VGND VGND VPWR VPWR U$$1096/Y sky130_fd_sc_hd__inv_1
XFILLER_149_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_81_7 U$$4026/X U$$4159/X U$$4292/X VGND VGND VPWR VPWR dadda_fa_2_82_3/B
+ dadda_fa_3_81_0/A sky130_fd_sc_hd__fa_2
XFILLER_144_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_74_6 U$$4145/X U$$4278/X U$$4411/X VGND VGND VPWR VPWR dadda_fa_2_75_2/B
+ dadda_fa_2_74_5/B sky130_fd_sc_hd__fa_1
XFILLER_59_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_5 input220/X dadda_fa_1_67_5/B dadda_fa_1_67_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_68_2/A dadda_fa_2_67_5/A sky130_fd_sc_hd__fa_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4116_1763 VGND VGND VPWR VPWR U$$4116_1763/HI U$$4116/A1 sky130_fd_sc_hd__conb_1
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_62_4 U$$1727/X U$$1860/X U$$1993/X VGND VGND VPWR VPWR dadda_fa_1_63_6/CIN
+ dadda_fa_1_62_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_40_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3905 U$$3905/A U$$3949/B VGND VGND VPWR VPWR U$$3905/X sky130_fd_sc_hd__xor2_1
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3916 U$$4053/A1 U$$3916/A2 U$$3916/B1 U$$3916/B2 VGND VGND VPWR VPWR U$$3917/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_19_2 U$$843/X U$$976/X VGND VGND VPWR VPWR dadda_fa_4_20_1/B dadda_ha_3_19_2/SUM
+ sky130_fd_sc_hd__ha_1
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3927 U$$3927/A U$$3935/B VGND VGND VPWR VPWR U$$3927/X sky130_fd_sc_hd__xor2_1
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$260 final_adder.U$$260/A final_adder.U$$260/B VGND VGND VPWR VPWR
+ final_adder.U$$322/B sky130_fd_sc_hd__and2_1
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$110 U$$382/B1 U$$118/A2 U$$384/B1 U$$118/B2 VGND VGND VPWR VPWR U$$111/A sky130_fd_sc_hd__a22o_1
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3938 U$$4075/A1 U$$3840/X U$$4214/A1 U$$3841/X VGND VGND VPWR VPWR U$$3939/A sky130_fd_sc_hd__a22o_1
XFILLER_100_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_604_ _613_/CLK _604_/D VGND VGND VPWR VPWR _604_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3949 U$$3949/A U$$3949/B VGND VGND VPWR VPWR U$$3949/X sky130_fd_sc_hd__xor2_1
XFILLER_73_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$271 final_adder.U$$270/A final_adder.U$$157/X final_adder.U$$159/X
+ VGND VGND VPWR VPWR final_adder.U$$271/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$282 final_adder.U$$282/A final_adder.U$$282/B VGND VGND VPWR VPWR
+ final_adder.U$$332/A sky130_fd_sc_hd__and2_1
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$121 U$$121/A U$$129/B VGND VGND VPWR VPWR U$$121/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_32_2 dadda_fa_3_32_2/A dadda_fa_3_32_2/B dadda_fa_3_32_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_1/A dadda_fa_4_32_2/B sky130_fd_sc_hd__fa_2
XFILLER_166_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$293 final_adder.U$$292/A final_adder.U$$201/X final_adder.U$$203/X
+ VGND VGND VPWR VPWR final_adder.U$$293/X sky130_fd_sc_hd__a21o_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$132 U$$406/A1 U$$4/X U$$406/B1 U$$5/X VGND VGND VPWR VPWR U$$133/A sky130_fd_sc_hd__a22o_1
XFILLER_40_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$143 U$$143/A1 U$$181/A2 U$$8/A1 U$$181/B2 VGND VGND VPWR VPWR U$$144/A sky130_fd_sc_hd__a22o_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$154 U$$154/A U$$180/B VGND VGND VPWR VPWR U$$154/X sky130_fd_sc_hd__xor2_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_25_1 U$$1121/X U$$1254/X U$$1387/X VGND VGND VPWR VPWR dadda_fa_4_26_0/CIN
+ dadda_fa_4_25_2/A sky130_fd_sc_hd__fa_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$165 U$$28/A1 U$$175/A2 U$$30/A1 U$$175/B2 VGND VGND VPWR VPWR U$$166/A sky130_fd_sc_hd__a22o_1
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_535_ _535_/CLK _535_/D VGND VGND VPWR VPWR _535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$176 U$$176/A U$$190/B VGND VGND VPWR VPWR U$$176/X sky130_fd_sc_hd__xor2_1
XFILLER_60_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$187 U$$733/B1 U$$219/A2 U$$600/A1 U$$219/B2 VGND VGND VPWR VPWR U$$188/A sky130_fd_sc_hd__a22o_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$198 U$$198/A U$$226/B VGND VGND VPWR VPWR U$$198/X sky130_fd_sc_hd__xor2_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_18_0 U$$43/X U$$176/X U$$309/X VGND VGND VPWR VPWR dadda_fa_4_19_1/A dadda_fa_4_18_2/A
+ sky130_fd_sc_hd__fa_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_466_ _466_/CLK _466_/D VGND VGND VPWR VPWR _466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_397_ _613_/CLK _397_/D VGND VGND VPWR VPWR _397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1252 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1010 U$$2877/A VGND VGND VPWR VPWR U$$2843/B sky130_fd_sc_hd__buf_6
XFILLER_86_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1021 U$$2541/B VGND VGND VPWR VPWR U$$2517/B sky130_fd_sc_hd__buf_8
XFILLER_142_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1032 U$$2442/B VGND VGND VPWR VPWR U$$2436/B sky130_fd_sc_hd__buf_6
Xrepeater1043 U$$2309/B VGND VGND VPWR VPWR U$$2269/B sky130_fd_sc_hd__buf_8
Xrepeater1054 U$$2174/B VGND VGND VPWR VPWR U$$2186/B sky130_fd_sc_hd__buf_8
XFILLER_142_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1065 U$$1870/B VGND VGND VPWR VPWR U$$1820/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_84_5 dadda_fa_2_84_5/A dadda_fa_2_84_5/B dadda_fa_2_84_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_2/A dadda_fa_4_84_0/A sky130_fd_sc_hd__fa_2
Xrepeater1076 U$$1719/B VGND VGND VPWR VPWR U$$1711/B sky130_fd_sc_hd__buf_8
Xrepeater1087 U$$1588/B VGND VGND VPWR VPWR U$$1578/B sky130_fd_sc_hd__buf_6
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1098 U$$1479/B VGND VGND VPWR VPWR U$$1501/B sky130_fd_sc_hd__buf_12
Xdadda_fa_2_77_4 dadda_fa_2_77_4/A dadda_fa_2_77_4/B dadda_fa_2_77_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/CIN dadda_fa_3_77_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_100_3 U$$3665/X U$$3798/X U$$3931/X VGND VGND VPWR VPWR dadda_fa_3_101_2/B
+ dadda_fa_3_100_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3020_1745 VGND VGND VPWR VPWR U$$3020_1745/HI U$$3020/A1 sky130_fd_sc_hd__conb_1
XFILLER_211_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_114_1 dadda_fa_5_114_1/A dadda_fa_5_114_1/B dadda_fa_5_114_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_115_0/B dadda_fa_7_114_0/A sky130_fd_sc_hd__fa_1
XFILLER_176_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_107_0 dadda_fa_5_107_0/A dadda_fa_5_107_0/B dadda_fa_5_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_108_0/A dadda_fa_6_107_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_17 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_110_0_1867 VGND VGND VPWR VPWR dadda_fa_3_110_0/A dadda_fa_3_110_0_1867/LO
+ sky130_fd_sc_hd__conb_1
Xdadda_fa_1_72_3 U$$3210/X U$$3343/X U$$3476/X VGND VGND VPWR VPWR dadda_fa_2_73_1/B
+ dadda_fa_2_72_4/B sky130_fd_sc_hd__fa_1
XFILLER_113_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_65_2 U$$3329/X U$$3462/X U$$3595/X VGND VGND VPWR VPWR dadda_fa_2_66_1/A
+ dadda_fa_2_65_4/A sky130_fd_sc_hd__fa_1
XFILLER_59_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_42_1 dadda_fa_4_42_1/A dadda_fa_4_42_1/B dadda_fa_4_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/B dadda_fa_5_42_1/B sky130_fd_sc_hd__fa_1
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_1 U$$1985/X U$$2118/X U$$2251/X VGND VGND VPWR VPWR dadda_fa_2_59_0/CIN
+ dadda_fa_2_58_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_115_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_35_0 dadda_fa_4_35_0/A dadda_fa_4_35_0/B dadda_fa_4_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/A dadda_fa_5_35_1/A sky130_fd_sc_hd__fa_1
XFILLER_55_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_320_ _442_/CLK _320_/D VGND VGND VPWR VPWR _320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_251_ _253_/CLK _251_/D VGND VGND VPWR VPWR _251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_182_ _189_/CLK _182_/D VGND VGND VPWR VPWR _182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_87_3 dadda_fa_3_87_3/A dadda_fa_3_87_3/B dadda_fa_3_87_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_1/B dadda_fa_4_87_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4403 U$$4403/A U$$4403/B VGND VGND VPWR VPWR U$$4403/X sky130_fd_sc_hd__xor2_1
XU$$4414 _563_/Q U$$4388/X U$$4416/A1 U$$4430/B2 VGND VGND VPWR VPWR U$$4415/A sky130_fd_sc_hd__a22o_1
XFILLER_38_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4425 U$$4425/A U$$4425/B VGND VGND VPWR VPWR U$$4425/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_60_1 U$$526/X U$$659/X U$$792/X VGND VGND VPWR VPWR dadda_fa_1_61_6/B
+ dadda_fa_1_60_8/A sky130_fd_sc_hd__fa_1
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4436 U$$4436/A1 U$$4388/X U$$4436/B1 U$$4496/B2 VGND VGND VPWR VPWR U$$4437/A
+ sky130_fd_sc_hd__a22o_1
XU$$4447 U$$4447/A U$$4447/B VGND VGND VPWR VPWR U$$4447/X sky130_fd_sc_hd__xor2_1
XFILLER_77_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3702 U$$3835/A U$$3702/B VGND VGND VPWR VPWR U$$3702/X sky130_fd_sc_hd__and2_1
XU$$4458 _585_/Q U$$4388/X _586_/Q U$$4468/B2 VGND VGND VPWR VPWR U$$4459/A sky130_fd_sc_hd__a22o_1
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3713 U$$3713/A1 U$$3743/A2 U$$3713/B1 U$$3743/B2 VGND VGND VPWR VPWR U$$3714/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3724 U$$3724/A U$$3832/B VGND VGND VPWR VPWR U$$3724/X sky130_fd_sc_hd__xor2_1
XU$$4469 U$$4469/A U$$4469/B VGND VGND VPWR VPWR U$$4469/X sky130_fd_sc_hd__xor2_1
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3735 U$$3735/A1 U$$3769/A2 U$$3735/B1 U$$3769/B2 VGND VGND VPWR VPWR U$$3736/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3746 U$$3746/A U$$3760/B VGND VGND VPWR VPWR U$$3746/X sky130_fd_sc_hd__xor2_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3757 _577_/Q U$$3785/A2 _578_/Q U$$3785/B2 VGND VGND VPWR VPWR U$$3758/A sky130_fd_sc_hd__a22o_1
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_109_2 dadda_fa_4_109_2/A dadda_fa_4_109_2/B dadda_fa_4_109_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/CIN dadda_fa_5_109_1/CIN sky130_fd_sc_hd__fa_1
XU$$3768 U$$3768/A U$$3816/B VGND VGND VPWR VPWR U$$3768/X sky130_fd_sc_hd__xor2_1
XU$$3779 U$$4464/A1 U$$3795/A2 U$$3779/B1 U$$3795/B2 VGND VGND VPWR VPWR U$$3780/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 U$$4176/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_361 U$$2812/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_518_ _520_/CLK _518_/D VGND VGND VPWR VPWR _518_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_372 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_383 _642_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_449_ _451_/CLK _449_/D VGND VGND VPWR VPWR _449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_82_2 dadda_fa_2_82_2/A dadda_fa_2_82_2/B dadda_fa_2_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/A dadda_fa_3_82_3/A sky130_fd_sc_hd__fa_1
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_75_1 dadda_fa_2_75_1/A dadda_fa_2_75_1/B dadda_fa_2_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_0/CIN dadda_fa_3_75_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_52_0 dadda_fa_5_52_0/A dadda_fa_5_52_0/B dadda_fa_5_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_53_0/A dadda_fa_6_52_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_68_0 dadda_fa_2_68_0/A dadda_fa_2_68_0/B dadda_fa_2_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_0/B dadda_fa_3_68_2/B sky130_fd_sc_hd__fa_1
XFILLER_69_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_97_2 dadda_fa_4_97_2/A dadda_fa_4_97_2/B dadda_fa_4_97_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/CIN dadda_fa_5_97_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_67_0 dadda_fa_7_67_0/A dadda_fa_7_67_0/B dadda_fa_7_67_0/CIN VGND VGND
+ VPWR VPWR _492_/D _363_/D sky130_fd_sc_hd__fa_1
XFILLER_191_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_70_0 U$$2275/X U$$2408/X U$$2541/X VGND VGND VPWR VPWR dadda_fa_2_71_0/B
+ dadda_fa_2_70_3/B sky130_fd_sc_hd__fa_1
XFILLER_132_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3009 U$$3283/A1 U$$2881/X U$$3285/A1 U$$2882/X VGND VGND VPWR VPWR U$$3010/A sky130_fd_sc_hd__a22o_1
XFILLER_75_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2308 U$$4361/B1 U$$2318/A2 U$$940/A1 U$$2318/B2 VGND VGND VPWR VPWR U$$2309/A
+ sky130_fd_sc_hd__a22o_1
XU$$2319 U$$2319/A U$$2321/B VGND VGND VPWR VPWR U$$2319/X sky130_fd_sc_hd__xor2_1
XFILLER_131_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1607 U$$922/A1 U$$1607/A2 U$$924/A1 U$$1607/B2 VGND VGND VPWR VPWR U$$1608/A sky130_fd_sc_hd__a22o_1
XU$$1618 U$$1618/A U$$1628/B VGND VGND VPWR VPWR U$$1618/X sky130_fd_sc_hd__xor2_1
XU$$1629 U$$2586/B1 U$$1635/A2 U$$2588/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1630/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk _628_/CLK VGND VGND VPWR VPWR _538_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_303_ _431_/CLK _303_/D VGND VGND VPWR VPWR _303_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_234_ _234_/CLK _234_/D VGND VGND VPWR VPWR _234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_92_1 dadda_fa_3_92_1/A dadda_fa_3_92_1/B dadda_fa_3_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_0/CIN dadda_fa_4_92_2/A sky130_fd_sc_hd__fa_1
XFILLER_109_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1069 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_85_0 dadda_fa_3_85_0/A dadda_fa_3_85_0/B dadda_fa_3_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_0/B dadda_fa_4_85_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_527 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater507 U$$3132/A2 VGND VGND VPWR VPWR U$$3120/A2 sky130_fd_sc_hd__buf_6
XFILLER_133_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater518 U$$2881/X VGND VGND VPWR VPWR U$$2973/A2 sky130_fd_sc_hd__buf_6
XFILLER_77_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4200 U$$4472/B1 U$$4202/A2 U$$4337/B1 U$$4202/B2 VGND VGND VPWR VPWR U$$4201/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater529 U$$2798/A2 VGND VGND VPWR VPWR U$$2788/A2 sky130_fd_sc_hd__buf_4
XFILLER_65_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4211 U$$4211/A U$$4247/A VGND VGND VPWR VPWR U$$4211/X sky130_fd_sc_hd__xor2_1
XU$$4222 U$$4222/A1 U$$4238/A2 U$$4498/A1 U$$4238/B2 VGND VGND VPWR VPWR U$$4223/A
+ sky130_fd_sc_hd__a22o_1
XU$$4233 U$$4233/A U$$4239/B VGND VGND VPWR VPWR U$$4233/X sky130_fd_sc_hd__xor2_1
XFILLER_120_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4244 U$$4516/B1 U$$4244/A2 U$$4244/B1 U$$4244/B2 VGND VGND VPWR VPWR U$$4245/A
+ sky130_fd_sc_hd__a22o_1
XU$$3510 U$$3510/A U$$3562/A VGND VGND VPWR VPWR U$$3510/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_114_0 U$$4092/X U$$4225/X U$$4358/X VGND VGND VPWR VPWR dadda_fa_5_115_0/A
+ dadda_fa_5_114_1/A sky130_fd_sc_hd__fa_1
XU$$4255 U$$4392/A1 U$$4297/A2 U$$4394/A1 U$$4297/B2 VGND VGND VPWR VPWR U$$4256/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_47_5 dadda_fa_2_47_5/A dadda_fa_2_47_5/B dadda_fa_2_47_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_2/A dadda_fa_4_47_0/A sky130_fd_sc_hd__fa_2
XU$$3521 U$$3658/A1 U$$3531/A2 U$$3521/B1 U$$3531/B2 VGND VGND VPWR VPWR U$$3522/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4266 U$$4266/A U$$4348/B VGND VGND VPWR VPWR U$$4266/X sky130_fd_sc_hd__xor2_1
XU$$4277 _563_/Q U$$4311/A2 U$$4416/A1 U$$4311/B2 VGND VGND VPWR VPWR U$$4278/A sky130_fd_sc_hd__a22o_1
XU$$3532 U$$3532/A U$$3538/B VGND VGND VPWR VPWR U$$3532/X sky130_fd_sc_hd__xor2_1
XFILLER_53_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4288 U$$4288/A U$$4296/B VGND VGND VPWR VPWR U$$4288/X sky130_fd_sc_hd__xor2_1
XU$$3543 U$$3952/B1 U$$3555/A2 U$$4228/B1 U$$3555/B2 VGND VGND VPWR VPWR U$$3544/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3554 U$$3554/A U$$3556/B VGND VGND VPWR VPWR U$$3554/X sky130_fd_sc_hd__xor2_1
XFILLER_80_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2820 U$$2957/A1 U$$2856/A2 U$$3916/B1 U$$2856/B2 VGND VGND VPWR VPWR U$$2821/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4299 _574_/Q U$$4347/A2 _575_/Q U$$4347/B2 VGND VGND VPWR VPWR U$$4300/A sky130_fd_sc_hd__a22o_1
XFILLER_80_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3565 _669_/Q U$$3565/B VGND VGND VPWR VPWR U$$3565/X sky130_fd_sc_hd__and2_1
XU$$3576 U$$3713/A1 U$$3612/A2 U$$3578/A1 U$$3612/B2 VGND VGND VPWR VPWR U$$3577/A
+ sky130_fd_sc_hd__a22o_1
XU$$2831 U$$2831/A U$$2843/B VGND VGND VPWR VPWR U$$2831/X sky130_fd_sc_hd__xor2_1
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3587 U$$3587/A U$$3609/B VGND VGND VPWR VPWR U$$3587/X sky130_fd_sc_hd__xor2_1
XU$$2842 U$$4075/A1 U$$2874/A2 U$$4214/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2843/A
+ sky130_fd_sc_hd__a22o_1
XU$$2853 U$$2853/A U$$2861/B VGND VGND VPWR VPWR U$$2853/X sky130_fd_sc_hd__xor2_1
XU$$3598 U$$3735/A1 U$$3636/A2 U$$3735/B1 U$$3636/B2 VGND VGND VPWR VPWR U$$3599/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2864 U$$2999/B1 U$$2866/A2 U$$2866/A1 U$$2866/B2 VGND VGND VPWR VPWR U$$2865/A
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_72_clk _634_/CLK VGND VGND VPWR VPWR _552_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_178_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2875 U$$2875/A U$$2875/B VGND VGND VPWR VPWR U$$2875/X sky130_fd_sc_hd__xor2_1
XU$$2886 U$$2886/A U$$2928/B VGND VGND VPWR VPWR U$$2886/X sky130_fd_sc_hd__xor2_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2897 U$$3445/A1 U$$2915/A2 U$$3310/A1 U$$2915/B2 VGND VGND VPWR VPWR U$$2898/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_180 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_1_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_33_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$709 U$$981/B1 U$$765/A2 U$$848/A1 U$$765/B2 VGND VGND VPWR VPWR U$$710/A sky130_fd_sc_hd__a22o_1
XFILLER_186_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_63_clk _535_/CLK VGND VGND VPWR VPWR _566_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1609 U$$4416/A1 VGND VGND VPWR VPWR U$$2909/A1 sky130_fd_sc_hd__buf_4
XFILLER_180_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_109_1 U$$3550/X U$$3683/X U$$3816/X VGND VGND VPWR VPWR dadda_fa_4_110_0/CIN
+ dadda_fa_4_109_2/A sky130_fd_sc_hd__fa_1
XFILLER_134_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1083 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2105 U$$3884/B1 U$$2109/A2 U$$3751/A1 U$$2109/B2 VGND VGND VPWR VPWR U$$2106/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2116 U$$2116/A U$$2144/B VGND VGND VPWR VPWR U$$2116/X sky130_fd_sc_hd__xor2_1
XU$$2127 U$$757/A1 U$$2135/A2 U$$759/A1 U$$2135/B2 VGND VGND VPWR VPWR U$$2128/A sky130_fd_sc_hd__a22o_1
XFILLER_90_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2138 U$$2138/A U$$2174/B VGND VGND VPWR VPWR U$$2138/X sky130_fd_sc_hd__xor2_1
XU$$1404 U$$2909/B1 U$$1442/A2 U$$2774/B1 U$$1442/B2 VGND VGND VPWR VPWR U$$1405/A
+ sky130_fd_sc_hd__a22o_1
XU$$2149 U$$916/A1 U$$2169/A2 U$$3519/B1 U$$2169/B2 VGND VGND VPWR VPWR U$$2150/A
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_54_clk _535_/CLK VGND VGND VPWR VPWR _526_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_27_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1415 U$$1415/A U$$1429/B VGND VGND VPWR VPWR U$$1415/X sky130_fd_sc_hd__xor2_1
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1426 U$$56/A1 U$$1458/A2 U$$467/B1 U$$1458/B2 VGND VGND VPWR VPWR U$$1427/A sky130_fd_sc_hd__a22o_1
XFILLER_188_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1437 U$$1437/A U$$1443/B VGND VGND VPWR VPWR U$$1437/X sky130_fd_sc_hd__xor2_1
XFILLER_203_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1448 U$$900/A1 U$$1486/A2 U$$4053/A1 U$$1486/B2 VGND VGND VPWR VPWR U$$1449/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1459 U$$1459/A U$$1459/B VGND VGND VPWR VPWR U$$1459/X sky130_fd_sc_hd__xor2_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_746 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_217_ _351_/CLK _217_/D VGND VGND VPWR VPWR _217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_52_3 dadda_fa_2_52_3/A dadda_fa_2_52_3/B dadda_fa_2_52_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/B dadda_fa_3_52_3/B sky130_fd_sc_hd__fa_1
XU$$4030 U$$4030/A U$$4044/B VGND VGND VPWR VPWR U$$4030/X sky130_fd_sc_hd__xor2_1
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4041 U$$4176/B1 U$$4071/A2 U$$4180/A1 U$$4071/B2 VGND VGND VPWR VPWR U$$4042/A
+ sky130_fd_sc_hd__a22o_1
XU$$4052 U$$4052/A U$$4058/B VGND VGND VPWR VPWR U$$4052/X sky130_fd_sc_hd__xor2_1
XFILLER_211_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4063 U$$4198/B1 U$$4071/A2 U$$4337/B1 U$$4071/B2 VGND VGND VPWR VPWR U$$4064/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_45_2 input196/X dadda_fa_2_45_2/B dadda_fa_2_45_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_46_1/A dadda_fa_3_45_3/A sky130_fd_sc_hd__fa_1
XFILLER_4_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4074 U$$4074/A U$$4084/B VGND VGND VPWR VPWR U$$4074/X sky130_fd_sc_hd__xor2_1
XU$$4085 U$$4222/A1 U$$4107/A2 U$$4087/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4086/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3340 U$$4160/B1 U$$3378/A2 U$$4027/A1 U$$3378/B2 VGND VGND VPWR VPWR U$$3341/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_22_1 dadda_fa_5_22_1/A dadda_fa_5_22_1/B dadda_fa_5_22_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_23_0/B dadda_fa_7_22_0/A sky130_fd_sc_hd__fa_1
XU$$3351 U$$3351/A U$$3357/B VGND VGND VPWR VPWR U$$3351/X sky130_fd_sc_hd__xor2_1
XU$$4096 U$$4096/A U$$4096/B VGND VGND VPWR VPWR U$$4096/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_38_1 U$$1546/X U$$1679/X U$$1812/X VGND VGND VPWR VPWR dadda_fa_3_39_0/CIN
+ dadda_fa_3_38_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_20_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3362 U$$3362/A1 U$$3378/A2 U$$3362/B1 U$$3378/B2 VGND VGND VPWR VPWR U$$3363/A
+ sky130_fd_sc_hd__a22o_1
XU$$3373 U$$3373/A U$$3424/A VGND VGND VPWR VPWR U$$3373/X sky130_fd_sc_hd__xor2_1
XU$$3384 U$$3658/A1 U$$3404/A2 U$$3521/B1 U$$3404/B2 VGND VGND VPWR VPWR U$$3385/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_45_clk _369_/CLK VGND VGND VPWR VPWR _504_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_202_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_15_0 dadda_fa_5_15_0/A dadda_fa_5_15_0/B dadda_fa_5_15_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_16_0/A dadda_fa_6_15_0/CIN sky130_fd_sc_hd__fa_1
XU$$3395 U$$3395/A U$$3397/B VGND VGND VPWR VPWR U$$3395/X sky130_fd_sc_hd__xor2_1
XU$$2650 U$$2650/A U$$2654/B VGND VGND VPWR VPWR U$$2650/X sky130_fd_sc_hd__xor2_1
XFILLER_206_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2661 U$$2796/B1 U$$2663/A2 U$$4168/B1 U$$2663/B2 VGND VGND VPWR VPWR U$$2662/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2672 U$$2672/A U$$2708/B VGND VGND VPWR VPWR U$$2672/X sky130_fd_sc_hd__xor2_1
XU$$2683 U$$2957/A1 U$$2687/A2 U$$3916/B1 U$$2687/B2 VGND VGND VPWR VPWR U$$2684/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2694 U$$2694/A U$$2734/B VGND VGND VPWR VPWR U$$2694/X sky130_fd_sc_hd__xor2_1
XFILLER_210_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1960 U$$999/B1 U$$2010/A2 U$$866/A1 U$$2010/B2 VGND VGND VPWR VPWR U$$1961/A sky130_fd_sc_hd__a22o_1
XFILLER_146_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1971 U$$1971/A U$$1977/B VGND VGND VPWR VPWR U$$1971/X sky130_fd_sc_hd__xor2_1
XFILLER_210_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1982 U$$749/A1 U$$1982/A2 U$$749/B1 U$$1982/B2 VGND VGND VPWR VPWR U$$1983/A sky130_fd_sc_hd__a22o_1
XFILLER_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1993 U$$1993/A U$$2003/B VGND VGND VPWR VPWR U$$1993/X sky130_fd_sc_hd__xor2_1
XFILLER_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput107 b[48] VGND VGND VPWR VPWR _600_/D sky130_fd_sc_hd__clkbuf_1
Xdadda_ha_1_41_3 U$$1286/X U$$1419/X VGND VGND VPWR VPWR dadda_fa_2_42_4/B dadda_fa_3_41_0/A
+ sky130_fd_sc_hd__ha_2
Xinput118 b[58] VGND VGND VPWR VPWR _610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput129 c[0] VGND VGND VPWR VPWR _424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_193_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$601 final_adder.U$$728/A final_adder.U$$728/B final_adder.U$$601/B1
+ VGND VGND VPWR VPWR final_adder.U$$729/B sky130_fd_sc_hd__a21o_1
XTAP_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1070 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$623 final_adder.U$$623/A final_adder.U$$623/B VGND VGND VPWR VPWR
+ _169_/D sky130_fd_sc_hd__xor2_1
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_4_11_1 U$$428/X U$$561/X VGND VGND VPWR VPWR dadda_fa_5_12_0/CIN dadda_ha_4_11_1/SUM
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$634 final_adder.U$$634/A final_adder.U$$634/B VGND VGND VPWR VPWR
+ _180_/D sky130_fd_sc_hd__xor2_4
XFILLER_186_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$645 final_adder.U$$645/A final_adder.U$$645/B VGND VGND VPWR VPWR
+ _191_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$656 final_adder.U$$656/A final_adder.U$$656/B VGND VGND VPWR VPWR
+ _202_/D sky130_fd_sc_hd__xor2_1
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater860 U$$217/B2 VGND VGND VPWR VPWR U$$249/B2 sky130_fd_sc_hd__buf_6
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$506 U$$506/A U$$518/B VGND VGND VPWR VPWR U$$506/X sky130_fd_sc_hd__xor2_1
Xrepeater871 U$$1375/X VGND VGND VPWR VPWR U$$1474/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$667 final_adder.U$$667/A final_adder.U$$667/B VGND VGND VPWR VPWR
+ _213_/D sky130_fd_sc_hd__xor2_4
XFILLER_99_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$678 final_adder.U$$678/A final_adder.U$$678/B VGND VGND VPWR VPWR
+ _224_/D sky130_fd_sc_hd__xor2_1
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$517 U$$791/A1 U$$517/A2 U$$517/B1 U$$517/B2 VGND VGND VPWR VPWR U$$518/A sky130_fd_sc_hd__a22o_1
Xrepeater882 U$$1190/B2 VGND VGND VPWR VPWR U$$1176/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_40_1 U$$486/X U$$619/X U$$752/X VGND VGND VPWR VPWR dadda_fa_2_41_4/A
+ dadda_fa_2_40_5/B sky130_fd_sc_hd__fa_1
XU$$528 U$$528/A U$$536/B VGND VGND VPWR VPWR U$$528/X sky130_fd_sc_hd__xor2_1
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater893 U$$98/B2 VGND VGND VPWR VPWR U$$128/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$689 final_adder.U$$689/A final_adder.U$$689/B VGND VGND VPWR VPWR
+ _235_/D sky130_fd_sc_hd__xor2_4
XFILLER_186_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$539 U$$676/A1 U$$545/A2 U$$676/B1 U$$545/B2 VGND VGND VPWR VPWR U$$540/A sky130_fd_sc_hd__a22o_1
XFILLER_71_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_clk _479_/CLK VGND VGND VPWR VPWR _353_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_80 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_91 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1406 U$$3916/B1 VGND VGND VPWR VPWR U$$3096/A1 sky130_fd_sc_hd__buf_6
Xrepeater1417 _588_/Q VGND VGND VPWR VPWR U$$4464/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1428 U$$896/B1 VGND VGND VPWR VPWR U$$76/A1 sky130_fd_sc_hd__buf_8
XFILLER_67_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1439 U$$4184/A1 VGND VGND VPWR VPWR U$$3088/A1 sky130_fd_sc_hd__buf_8
XFILLER_106_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_62_2 dadda_fa_3_62_2/A dadda_fa_3_62_2/B dadda_fa_3_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_1/A dadda_fa_4_62_2/B sky130_fd_sc_hd__fa_1
XFILLER_79_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_55_1 dadda_fa_3_55_1/A dadda_fa_3_55_1/B dadda_fa_3_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_0/CIN dadda_fa_4_55_2/A sky130_fd_sc_hd__fa_1
XFILLER_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_32_0 dadda_fa_6_32_0/A dadda_fa_6_32_0/B dadda_fa_6_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_33_0/B dadda_fa_7_32_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_36_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_48_0 dadda_fa_3_48_0/A dadda_fa_3_48_0/B dadda_fa_3_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_0/B dadda_fa_4_48_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_36_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk _432_/CLK VGND VGND VPWR VPWR _207_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_165_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1201 U$$1201/A U$$1203/B VGND VGND VPWR VPWR U$$1201/X sky130_fd_sc_hd__xor2_1
XFILLER_16_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1212 U$$2171/A1 U$$1230/A2 U$$392/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1213/A
+ sky130_fd_sc_hd__a22o_1
XU$$1223 U$$1223/A U$$1225/B VGND VGND VPWR VPWR U$$1223/X sky130_fd_sc_hd__xor2_1
XFILLER_16_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1234 _634_/Q VGND VGND VPWR VPWR U$$1236/B sky130_fd_sc_hd__inv_1
XFILLER_62_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1245 U$$12/A1 U$$1279/A2 U$$14/A1 U$$1279/B2 VGND VGND VPWR VPWR U$$1246/A sky130_fd_sc_hd__a22o_1
XU$$1256 U$$1256/A U$$1292/B VGND VGND VPWR VPWR U$$1256/X sky130_fd_sc_hd__xor2_1
XU$$1267 U$$582/A1 U$$1279/A2 U$$582/B1 U$$1279/B2 VGND VGND VPWR VPWR U$$1268/A sky130_fd_sc_hd__a22o_1
XU$$1278 U$$1278/A U$$1280/B VGND VGND VPWR VPWR U$$1278/X sky130_fd_sc_hd__xor2_1
XU$$1289 U$$330/A1 U$$1323/A2 U$$2796/B1 U$$1323/B2 VGND VGND VPWR VPWR U$$1290/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1046 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_105_0 dadda_fa_7_105_0/A dadda_fa_7_105_0/B dadda_fa_7_105_0/CIN VGND
+ VGND VPWR VPWR _530_/D _401_/D sky130_fd_sc_hd__fa_1
XFILLER_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_50_0 U$$3478/B input202/X dadda_fa_2_50_0/CIN VGND VGND VPWR VPWR dadda_fa_3_51_0/B
+ dadda_fa_3_50_2/B sky130_fd_sc_hd__fa_1
XFILLER_61_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3170 U$$3170/A U$$3218/B VGND VGND VPWR VPWR U$$3170/X sky130_fd_sc_hd__xor2_1
XU$$3181 U$$3453/B1 U$$3209/A2 U$$3181/B1 U$$3209/B2 VGND VGND VPWR VPWR U$$3182/A
+ sky130_fd_sc_hd__a22o_1
XU$$3192 U$$3192/A U$$3236/B VGND VGND VPWR VPWR U$$3192/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_94_0_1861 VGND VGND VPWR VPWR dadda_fa_1_94_0/A dadda_fa_1_94_0_1861/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_50_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2480 U$$562/A1 U$$2530/A2 U$$3713/B1 U$$2530/B2 VGND VGND VPWR VPWR U$$2481/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2491 U$$2491/A U$$2541/B VGND VGND VPWR VPWR U$$2491/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1790 U$$1790/A U$$1820/B VGND VGND VPWR VPWR U$$1790/X sky130_fd_sc_hd__xor2_1
XFILLER_22_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_72_1 dadda_fa_4_72_1/A dadda_fa_4_72_1/B dadda_fa_4_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/B dadda_fa_5_72_1/B sky130_fd_sc_hd__fa_1
XFILLER_116_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_88_1 U$$2045/X U$$2178/X U$$2311/X VGND VGND VPWR VPWR dadda_fa_2_89_3/CIN
+ dadda_fa_2_88_5/A sky130_fd_sc_hd__fa_1
XFILLER_150_549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_65_0 dadda_fa_4_65_0/A dadda_fa_4_65_0/B dadda_fa_4_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/A dadda_fa_5_65_1/A sky130_fd_sc_hd__fa_1
XFILLER_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_999 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_620_ _624_/CLK _620_/D VGND VGND VPWR VPWR _620_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$431 final_adder.U$$348/B final_adder.U$$734/B final_adder.U$$313/X
+ VGND VGND VPWR VPWR final_adder.U$$738/B sky130_fd_sc_hd__a21o_2
Xdadda_fa_0_68_0_1849 VGND VGND VPWR VPWR dadda_fa_0_68_0/A dadda_fa_0_68_0_1849/LO
+ sky130_fd_sc_hd__conb_1
XTAP_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$453 final_adder.U$$276/B final_adder.U$$662/B final_adder.U$$169/X
+ VGND VGND VPWR VPWR final_adder.U$$664/B sky130_fd_sc_hd__a21o_1
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$303 U$$303/A U$$335/B VGND VGND VPWR VPWR U$$303/X sky130_fd_sc_hd__xor2_1
XFILLER_45_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$475 final_adder.U$$298/B final_adder.U$$706/B final_adder.U$$213/X
+ VGND VGND VPWR VPWR final_adder.U$$708/B sky130_fd_sc_hd__a21o_1
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$314 U$$449/B1 U$$318/A2 U$$316/A1 U$$318/B2 VGND VGND VPWR VPWR U$$315/A sky130_fd_sc_hd__a22o_1
XFILLER_45_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$325 U$$325/A U$$335/B VGND VGND VPWR VPWR U$$325/X sky130_fd_sc_hd__xor2_1
X_551_ _627_/CLK _551_/D VGND VGND VPWR VPWR _551_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater690 U$$4115/X VGND VGND VPWR VPWR U$$4244/B2 sky130_fd_sc_hd__buf_4
XFILLER_205_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$497 final_adder.U$$624/A final_adder.U$$624/B final_adder.U$$497/B1
+ VGND VGND VPWR VPWR final_adder.U$$625/B sky130_fd_sc_hd__a21o_1
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$336 U$$882/B1 U$$350/A2 U$$747/B1 U$$350/B2 VGND VGND VPWR VPWR U$$337/A sky130_fd_sc_hd__a22o_1
XU$$347 U$$347/A U$$351/B VGND VGND VPWR VPWR U$$347/X sky130_fd_sc_hd__xor2_1
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$358 U$$358/A1 U$$398/A2 U$$86/A1 U$$398/B2 VGND VGND VPWR VPWR U$$359/A sky130_fd_sc_hd__a22o_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$369 U$$369/A U$$383/B VGND VGND VPWR VPWR U$$369/X sky130_fd_sc_hd__xor2_1
X_482_ _482_/CLK _482_/D VGND VGND VPWR VPWR _482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1046 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4501_1829 VGND VGND VPWR VPWR U$$4501_1829/HI U$$4501/B sky130_fd_sc_hd__conb_1
XFILLER_41_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1203 U$$2459/B1 VGND VGND VPWR VPWR U$$678/B1 sky130_fd_sc_hd__buf_6
XFILLER_165_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1214 _613_/Q VGND VGND VPWR VPWR U$$3281/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1225 U$$811/A1 VGND VGND VPWR VPWR U$$674/A1 sky130_fd_sc_hd__buf_6
Xrepeater1236 U$$3412/A1 VGND VGND VPWR VPWR U$$4369/B1 sky130_fd_sc_hd__buf_4
Xrepeater1247 _609_/Q VGND VGND VPWR VPWR U$$2725/A1 sky130_fd_sc_hd__buf_6
XFILLER_154_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1258 U$$4500/B1 VGND VGND VPWR VPWR U$$938/B1 sky130_fd_sc_hd__buf_6
XFILLER_181_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4393_1775 VGND VGND VPWR VPWR U$$4393_1775/HI U$$4393/B sky130_fd_sc_hd__conb_1
Xrepeater1269 U$$3404/A1 VGND VGND VPWR VPWR U$$4087/B1 sky130_fd_sc_hd__buf_6
XFILLER_136_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4469_1813 VGND VGND VPWR VPWR U$$4469_1813/HI U$$4469/B sky130_fd_sc_hd__conb_1
XFILLER_122_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_636 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_864 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$870 U$$48/A1 U$$878/A2 U$$48/B1 U$$878/B2 VGND VGND VPWR VPWR U$$871/A sky130_fd_sc_hd__a22o_1
XFILLER_91_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1020 U$$1020/A U$$996/B VGND VGND VPWR VPWR U$$1020/X sky130_fd_sc_hd__xor2_1
XFILLER_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$881 U$$881/A U$$897/B VGND VGND VPWR VPWR U$$881/X sky130_fd_sc_hd__xor2_1
XFILLER_211_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$892 U$$70/A1 U$$924/A2 U$$894/A1 U$$924/B2 VGND VGND VPWR VPWR U$$893/A sky130_fd_sc_hd__a22o_1
XFILLER_91_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1031 U$$894/A1 U$$1039/A2 U$$896/A1 U$$1039/B2 VGND VGND VPWR VPWR U$$1032/A sky130_fd_sc_hd__a22o_1
XU$$1042 U$$1042/A U$$1090/B VGND VGND VPWR VPWR U$$1042/X sky130_fd_sc_hd__xor2_1
XFILLER_50_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1053 U$$94/A1 U$$997/A2 U$$96/A1 U$$997/B2 VGND VGND VPWR VPWR U$$1054/A sky130_fd_sc_hd__a22o_1
XU$$1064 U$$1064/A U$$996/B VGND VGND VPWR VPWR U$$1064/X sky130_fd_sc_hd__xor2_1
XFILLER_56_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1075 U$$527/A1 U$$963/X U$$392/A1 U$$964/X VGND VGND VPWR VPWR U$$1076/A sky130_fd_sc_hd__a22o_1
XFILLER_91_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1086 U$$1086/A U$$1095/A VGND VGND VPWR VPWR U$$1086/X sky130_fd_sc_hd__xor2_1
XFILLER_148_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1097 _632_/Q VGND VGND VPWR VPWR U$$1099/B sky130_fd_sc_hd__inv_1
XFILLER_32_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1042 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_82_0 dadda_fa_5_82_0/A dadda_fa_5_82_0/B dadda_fa_5_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_83_0/A dadda_fa_6_82_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_144_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_98_0 dadda_fa_2_98_0/A U$$2464/X U$$2597/X VGND VGND VPWR VPWR dadda_fa_3_99_0/CIN
+ dadda_fa_3_98_2/B sky130_fd_sc_hd__fa_1
XFILLER_105_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_7_clk _442_/CLK VGND VGND VPWR VPWR _435_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_579 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_74_7 input228/X dadda_fa_1_74_7/B dadda_fa_1_74_7/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_75_2/CIN dadda_fa_2_74_5/CIN sky130_fd_sc_hd__fa_2
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_67_6 dadda_fa_1_67_6/A dadda_fa_1_67_6/B dadda_fa_1_67_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_2/B dadda_fa_2_67_5/B sky130_fd_sc_hd__fa_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1040 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_94_1 U$$2456/X U$$2589/X VGND VGND VPWR VPWR dadda_fa_2_95_5/CIN dadda_fa_3_94_0/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_7_97_0 dadda_fa_7_97_0/A dadda_fa_7_97_0/B dadda_fa_7_97_0/CIN VGND VGND
+ VPWR VPWR _522_/D _393_/D sky130_fd_sc_hd__fa_1
XFILLER_195_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1030 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_803 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_112_0 dadda_fa_6_112_0/A dadda_fa_6_112_0/B dadda_fa_6_112_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_113_0/B dadda_fa_7_112_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3906 U$$4180/A1 U$$3910/A2 U$$4045/A1 U$$3910/B2 VGND VGND VPWR VPWR U$$3907/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3917 U$$3917/A U$$3917/B VGND VGND VPWR VPWR U$$3917/X sky130_fd_sc_hd__xor2_1
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3928 _594_/Q U$$3932/A2 U$$4065/B1 U$$3932/B2 VGND VGND VPWR VPWR U$$3929/A sky130_fd_sc_hd__a22o_1
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$250 final_adder.U$$745/A final_adder.U$$744/A VGND VGND VPWR VPWR
+ final_adder.U$$316/A sky130_fd_sc_hd__and2_1
X_603_ _613_/CLK _603_/D VGND VGND VPWR VPWR _603_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$261 final_adder.U$$260/A final_adder.U$$137/X final_adder.U$$139/X
+ VGND VGND VPWR VPWR final_adder.U$$261/X sky130_fd_sc_hd__a21o_1
XU$$3939 U$$3939/A U$$3943/B VGND VGND VPWR VPWR U$$3939/X sky130_fd_sc_hd__xor2_1
XU$$100 U$$98/B1 U$$98/A2 U$$648/B1 U$$98/B2 VGND VGND VPWR VPWR U$$101/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$272 final_adder.U$$272/A final_adder.U$$272/B VGND VGND VPWR VPWR
+ final_adder.U$$328/B sky130_fd_sc_hd__and2_1
XU$$111 U$$111/A U$$117/B VGND VGND VPWR VPWR U$$111/X sky130_fd_sc_hd__xor2_1
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$283 final_adder.U$$282/A final_adder.U$$181/X final_adder.U$$183/X
+ VGND VGND VPWR VPWR final_adder.U$$283/X sky130_fd_sc_hd__a21o_1
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_32_3 dadda_fa_3_32_3/A dadda_fa_3_32_3/B dadda_fa_3_32_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_1/B dadda_fa_4_32_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$122 U$$942/B1 U$$128/A2 U$$946/A1 U$$128/B2 VGND VGND VPWR VPWR U$$123/A sky130_fd_sc_hd__a22o_1
XFILLER_206_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$294 final_adder.U$$294/A final_adder.U$$294/B VGND VGND VPWR VPWR
+ final_adder.U$$338/A sky130_fd_sc_hd__and2_1
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$133 U$$133/A U$$2/A VGND VGND VPWR VPWR U$$133/X sky130_fd_sc_hd__xor2_1
XU$$144 U$$144/A U$$180/B VGND VGND VPWR VPWR U$$144/X sky130_fd_sc_hd__xor2_1
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$155 U$$429/A1 U$$175/A2 U$$429/B1 U$$175/B2 VGND VGND VPWR VPWR U$$156/A sky130_fd_sc_hd__a22o_1
X_534_ _534_/CLK _534_/D VGND VGND VPWR VPWR _534_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$166 U$$166/A U$$190/B VGND VGND VPWR VPWR U$$166/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_25_2 U$$1520/X U$$1653/X input174/X VGND VGND VPWR VPWR dadda_fa_4_26_1/A
+ dadda_fa_4_25_2/B sky130_fd_sc_hd__fa_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$177 U$$449/B1 U$$181/A2 U$$316/A1 U$$181/B2 VGND VGND VPWR VPWR U$$178/A sky130_fd_sc_hd__a22o_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$188 U$$188/A U$$190/B VGND VGND VPWR VPWR U$$188/X sky130_fd_sc_hd__xor2_1
XU$$199 U$$62/A1 U$$219/A2 U$$64/A1 U$$219/B2 VGND VGND VPWR VPWR U$$200/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_18_1 U$$442/X U$$575/X U$$708/X VGND VGND VPWR VPWR dadda_fa_4_19_1/B
+ dadda_fa_4_18_2/B sky130_fd_sc_hd__fa_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_465_ _466_/CLK _465_/D VGND VGND VPWR VPWR _465_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4499_1828 VGND VGND VPWR VPWR U$$4499_1828/HI U$$4499/B sky130_fd_sc_hd__conb_1
XFILLER_129_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_396_ _613_/CLK _396_/D VGND VGND VPWR VPWR _396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_619 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1000 U$$2972/B VGND VGND VPWR VPWR U$$2928/B sky130_fd_sc_hd__buf_6
XFILLER_154_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1011 _657_/Q VGND VGND VPWR VPWR U$$2877/A sky130_fd_sc_hd__buf_6
XFILLER_126_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1022 U$$2567/B VGND VGND VPWR VPWR U$$2551/B sky130_fd_sc_hd__buf_6
XFILLER_5_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1033 U$$2388/B VGND VGND VPWR VPWR U$$2366/B sky130_fd_sc_hd__buf_8
XFILLER_99_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1044 U$$2321/B VGND VGND VPWR VPWR U$$2328/A sky130_fd_sc_hd__buf_6
XFILLER_5_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1055 _647_/Q VGND VGND VPWR VPWR U$$2174/B sky130_fd_sc_hd__buf_6
XFILLER_175_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1066 U$$1918/A VGND VGND VPWR VPWR U$$1870/B sky130_fd_sc_hd__buf_6
Xrepeater1077 U$$1747/B VGND VGND VPWR VPWR U$$1719/B sky130_fd_sc_hd__buf_6
XFILLER_142_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_590 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1088 U$$1588/B VGND VGND VPWR VPWR U$$1562/B sky130_fd_sc_hd__buf_6
Xrepeater1099 U$$1507/A VGND VGND VPWR VPWR U$$1479/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_77_5 dadda_fa_2_77_5/A dadda_fa_2_77_5/B dadda_fa_2_77_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_2/A dadda_fa_4_77_0/A sky130_fd_sc_hd__fa_2
XFILLER_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_107_1 dadda_fa_5_107_1/A dadda_fa_5_107_1/B dadda_fa_5_107_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_108_0/B dadda_fa_7_107_0/A sky130_fd_sc_hd__fa_2
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_72_4 U$$3609/X U$$3742/X U$$3875/X VGND VGND VPWR VPWR dadda_fa_2_73_1/CIN
+ dadda_fa_2_72_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_65_3 U$$3728/X U$$3861/X U$$3994/X VGND VGND VPWR VPWR dadda_fa_2_66_1/B
+ dadda_fa_2_65_4/B sky130_fd_sc_hd__fa_1
XFILLER_63_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_42_2 dadda_fa_4_42_2/A dadda_fa_4_42_2/B dadda_fa_4_42_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/CIN dadda_fa_5_42_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_2 U$$2384/X U$$2517/X U$$2650/X VGND VGND VPWR VPWR dadda_fa_2_59_1/A
+ dadda_fa_2_58_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_35_1 dadda_fa_4_35_1/A dadda_fa_4_35_1/B dadda_fa_4_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/B dadda_fa_5_35_1/B sky130_fd_sc_hd__fa_1
XFILLER_64_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_12_0 dadda_fa_7_12_0/A dadda_fa_7_12_0/B dadda_fa_7_12_0/CIN VGND VGND
+ VPWR VPWR _437_/D _308_/D sky130_fd_sc_hd__fa_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_28_0 dadda_fa_4_28_0/A dadda_fa_4_28_0/B dadda_fa_4_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/A dadda_fa_5_28_1/A sky130_fd_sc_hd__fa_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_250_ _253_/CLK _250_/D VGND VGND VPWR VPWR _250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_181_ _189_/CLK _181_/D VGND VGND VPWR VPWR _181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_0_61_4 U$$1725/X U$$1858/X VGND VGND VPWR VPWR dadda_fa_1_62_7/A dadda_fa_2_61_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_124_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4404 U$$4404/A1 U$$4388/X U$$4404/B1 U$$4430/B2 VGND VGND VPWR VPWR U$$4405/A
+ sky130_fd_sc_hd__a22o_1
XU$$4415 U$$4415/A U$$4415/B VGND VGND VPWR VPWR U$$4415/X sky130_fd_sc_hd__xor2_1
XFILLER_78_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_60_2 U$$925/X U$$1058/X U$$1191/X VGND VGND VPWR VPWR dadda_fa_1_61_6/CIN
+ dadda_fa_1_60_8/B sky130_fd_sc_hd__fa_1
XFILLER_65_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4426 U$$4426/A1 U$$4388/X _570_/Q U$$4454/B2 VGND VGND VPWR VPWR U$$4427/A sky130_fd_sc_hd__a22o_1
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4437 U$$4437/A U$$4437/B VGND VGND VPWR VPWR U$$4437/X sky130_fd_sc_hd__xor2_1
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3703 U$$3701/Y _670_/Q U$$3699/A U$$3702/X U$$3699/Y VGND VGND VPWR VPWR U$$3703/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_93_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4448 U$$4448/A1 U$$4388/X U$$4450/A1 U$$4454/B2 VGND VGND VPWR VPWR U$$4449/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4459 U$$4459/A U$$4459/B VGND VGND VPWR VPWR U$$4459/X sky130_fd_sc_hd__xor2_1
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3714 U$$3714/A U$$3764/B VGND VGND VPWR VPWR U$$3714/X sky130_fd_sc_hd__xor2_1
XFILLER_206_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3725 U$$4136/A1 U$$3833/A2 U$$4136/B1 U$$3833/B2 VGND VGND VPWR VPWR U$$3726/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3736 U$$3736/A U$$3816/B VGND VGND VPWR VPWR U$$3736/X sky130_fd_sc_hd__xor2_1
XU$$3747 U$$4156/B1 U$$3785/A2 U$$3884/B1 U$$3785/B2 VGND VGND VPWR VPWR U$$3748/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3758 U$$3758/A U$$3800/B VGND VGND VPWR VPWR U$$3758/X sky130_fd_sc_hd__xor2_1
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_0 U$$1929/X U$$2062/X U$$2130/B VGND VGND VPWR VPWR dadda_fa_4_31_0/B
+ dadda_fa_4_30_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_205_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_1011 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3769 U$$3769/A1 U$$3769/A2 U$$3769/B1 U$$3769/B2 VGND VGND VPWR VPWR U$$3770/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_340 U$$3112/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_351 U$$749/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_517_ _520_/CLK _517_/D VGND VGND VPWR VPWR _517_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_362 U$$2040/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1028 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_373 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_384 _644_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_448_ _448_/CLK _448_/D VGND VGND VPWR VPWR _448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_379_ _379_/CLK _379_/D VGND VGND VPWR VPWR _379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_983 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_82_3 dadda_fa_2_82_3/A dadda_fa_2_82_3/B dadda_fa_2_82_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/B dadda_fa_3_82_3/B sky130_fd_sc_hd__fa_1
XFILLER_170_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_75_2 dadda_fa_2_75_2/A dadda_fa_2_75_2/B dadda_fa_2_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/A dadda_fa_3_75_3/A sky130_fd_sc_hd__fa_1
XFILLER_141_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_52_1 dadda_fa_5_52_1/A dadda_fa_5_52_1/B dadda_fa_5_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_53_0/B dadda_fa_7_52_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_68_1 dadda_fa_2_68_1/A dadda_fa_2_68_1/B dadda_fa_2_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_0/CIN dadda_fa_3_68_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_45_0 dadda_fa_5_45_0/A dadda_fa_5_45_0/B dadda_fa_5_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_46_0/A dadda_fa_6_45_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_70_1 U$$2674/X U$$2807/X U$$2940/X VGND VGND VPWR VPWR dadda_fa_2_71_0/CIN
+ dadda_fa_2_70_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1056 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_63_0 U$$2394/X U$$2527/X U$$2660/X VGND VGND VPWR VPWR dadda_fa_2_64_0/B
+ dadda_fa_2_63_3/B sky130_fd_sc_hd__fa_1
XFILLER_75_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2309 U$$2309/A U$$2309/B VGND VGND VPWR VPWR U$$2309/X sky130_fd_sc_hd__xor2_1
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1608 U$$1608/A U$$1642/B VGND VGND VPWR VPWR U$$1608/X sky130_fd_sc_hd__xor2_1
XU$$1619 U$$3124/B1 U$$1627/A2 U$$2991/A1 U$$1627/B2 VGND VGND VPWR VPWR U$$1620/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_131_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_302_ _428_/CLK _302_/D VGND VGND VPWR VPWR _302_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_233_ _234_/CLK _233_/D VGND VGND VPWR VPWR _233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_92_2 dadda_fa_3_92_2/A dadda_fa_3_92_2/B dadda_fa_3_92_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_1/A dadda_fa_4_92_2/B sky130_fd_sc_hd__fa_1
XFILLER_108_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_85_1 dadda_fa_3_85_1/A dadda_fa_3_85_1/B dadda_fa_3_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_0/CIN dadda_fa_4_85_2/A sky130_fd_sc_hd__fa_1
XFILLER_124_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_62_0 dadda_fa_6_62_0/A dadda_fa_6_62_0/B dadda_fa_6_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_63_0/B dadda_fa_7_62_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_78_0 dadda_fa_3_78_0/A dadda_fa_3_78_0/B dadda_fa_3_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_0/B dadda_fa_4_78_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_ha_0_52_0 U$$111/X U$$244/X VGND VGND VPWR VPWR dadda_fa_1_53_8/CIN dadda_fa_2_52_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_97_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater508 U$$3144/A2 VGND VGND VPWR VPWR U$$3132/A2 sky130_fd_sc_hd__buf_4
XU$$4201 U$$4201/A U$$4203/B VGND VGND VPWR VPWR U$$4201/X sky130_fd_sc_hd__xor2_1
Xrepeater519 U$$308/A2 VGND VGND VPWR VPWR U$$318/A2 sky130_fd_sc_hd__buf_4
XU$$4212 U$$4486/A1 U$$4244/A2 U$$4351/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4213/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4223 U$$4223/A U$$4246/A VGND VGND VPWR VPWR U$$4223/X sky130_fd_sc_hd__xor2_1
XU$$4234 U$$4369/B1 U$$4238/A2 U$$4236/A1 U$$4238/B2 VGND VGND VPWR VPWR U$$4235/A
+ sky130_fd_sc_hd__a22o_1
XU$$4245 U$$4245/A U$$4246/A VGND VGND VPWR VPWR U$$4245/X sky130_fd_sc_hd__xor2_1
XU$$3500 U$$3500/A U$$3506/B VGND VGND VPWR VPWR U$$3500/X sky130_fd_sc_hd__xor2_1
XU$$4256 U$$4256/A U$$4298/B VGND VGND VPWR VPWR U$$4256/X sky130_fd_sc_hd__xor2_1
XU$$3511 U$$4470/A1 U$$3429/X U$$4333/B1 U$$3430/X VGND VGND VPWR VPWR U$$3512/A sky130_fd_sc_hd__a22o_1
XU$$3522 U$$3522/A U$$3538/B VGND VGND VPWR VPWR U$$3522/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_114_1 U$$4491/X input145/X dadda_fa_4_114_1/CIN VGND VGND VPWR VPWR dadda_fa_5_115_0/B
+ dadda_fa_5_114_1/B sky130_fd_sc_hd__fa_1
XU$$4267 _558_/Q U$$4297/A2 U$$4404/B1 U$$4297/B2 VGND VGND VPWR VPWR U$$4268/A sky130_fd_sc_hd__a22o_1
XFILLER_20_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4278 U$$4278/A U$$4296/B VGND VGND VPWR VPWR U$$4278/X sky130_fd_sc_hd__xor2_1
XU$$3533 U$$3805/B1 U$$3537/A2 U$$3807/B1 U$$3537/B2 VGND VGND VPWR VPWR U$$3534/A
+ sky130_fd_sc_hd__a22o_1
XU$$4289 _569_/Q U$$4311/A2 _570_/Q U$$4311/B2 VGND VGND VPWR VPWR U$$4290/A sky130_fd_sc_hd__a22o_1
XU$$3544 U$$3544/A U$$3556/B VGND VGND VPWR VPWR U$$3544/X sky130_fd_sc_hd__xor2_1
XU$$3555 U$$4514/A1 U$$3555/A2 U$$4516/A1 U$$3555/B2 VGND VGND VPWR VPWR U$$3556/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2810 U$$3495/A1 U$$2812/A2 U$$4317/B1 U$$2812/B2 VGND VGND VPWR VPWR U$$2811/A
+ sky130_fd_sc_hd__a22o_1
XU$$2821 U$$2821/A U$$2861/B VGND VGND VPWR VPWR U$$2821/X sky130_fd_sc_hd__xor2_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_107_0 dadda_fa_4_107_0/A dadda_fa_4_107_0/B dadda_fa_4_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/A dadda_fa_5_107_1/A sky130_fd_sc_hd__fa_1
XU$$3566 U$$3564/Y _668_/Q _667_/Q U$$3565/X U$$3562/Y VGND VGND VPWR VPWR U$$3566/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_92_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3577 U$$3577/A U$$3613/B VGND VGND VPWR VPWR U$$3577/X sky130_fd_sc_hd__xor2_1
XFILLER_19_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2832 U$$3380/A1 U$$2832/A2 U$$2832/B1 U$$2832/B2 VGND VGND VPWR VPWR U$$2833/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2843 U$$2843/A U$$2843/B VGND VGND VPWR VPWR U$$2843/X sky130_fd_sc_hd__xor2_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3588 U$$4136/A1 U$$3628/A2 U$$4136/B1 U$$3628/B2 VGND VGND VPWR VPWR U$$3589/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2854 U$$2991/A1 U$$2856/A2 U$$2991/B1 U$$2856/B2 VGND VGND VPWR VPWR U$$2855/A
+ sky130_fd_sc_hd__a22o_1
XU$$3599 U$$3599/A U$$3637/B VGND VGND VPWR VPWR U$$3599/X sky130_fd_sc_hd__xor2_1
XU$$2865 U$$2865/A _657_/Q VGND VGND VPWR VPWR U$$2865/X sky130_fd_sc_hd__xor2_1
XFILLER_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2876 U$$2877/A VGND VGND VPWR VPWR U$$2876/Y sky130_fd_sc_hd__inv_1
XFILLER_209_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_170 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2887 U$$3022/B1 U$$2929/A2 U$$3024/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2888/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2898 U$$2898/A U$$2916/B VGND VGND VPWR VPWR U$$2898/X sky130_fd_sc_hd__xor2_1
XFILLER_60_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_181 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_80_0 input235/X dadda_fa_2_80_0/B dadda_fa_2_80_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_81_0/B dadda_fa_3_80_2/B sky130_fd_sc_hd__fa_1
XFILLER_88_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_50_8 U$$3299/X U$$3432/X VGND VGND VPWR VPWR dadda_fa_2_51_3/A dadda_fa_3_50_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_142_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$143_1719 VGND VGND VPWR VPWR U$$143_1719/HI U$$143/A1 sky130_fd_sc_hd__conb_1
XFILLER_71_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_95_0 dadda_fa_4_95_0/A dadda_fa_4_95_0/B dadda_fa_4_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/A dadda_fa_5_95_1/A sky130_fd_sc_hd__fa_1
XFILLER_193_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_109_2 U$$3949/X U$$4082/X U$$4215/X VGND VGND VPWR VPWR dadda_fa_4_110_1/A
+ dadda_fa_4_109_2/B sky130_fd_sc_hd__fa_1
XFILLER_69_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput380 _264_/Q VGND VGND VPWR VPWR o[96] sky130_fd_sc_hd__buf_2
XFILLER_43_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2106 U$$2106/A U$$2108/B VGND VGND VPWR VPWR U$$2106/X sky130_fd_sc_hd__xor2_1
XFILLER_75_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2117 U$$334/B1 U$$2145/A2 U$$201/A1 U$$2145/B2 VGND VGND VPWR VPWR U$$2118/A sky130_fd_sc_hd__a22o_1
XFILLER_16_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2128 U$$2128/A U$$2136/B VGND VGND VPWR VPWR U$$2128/X sky130_fd_sc_hd__xor2_1
XFILLER_76_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2139 U$$3372/A1 U$$2059/X U$$3374/A1 U$$2060/X VGND VGND VPWR VPWR U$$2140/A sky130_fd_sc_hd__a22o_1
XFILLER_90_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1405 U$$1405/A U$$1443/B VGND VGND VPWR VPWR U$$1405/X sky130_fd_sc_hd__xor2_1
XFILLER_167_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1416 U$$729/B1 U$$1424/A2 U$$733/A1 U$$1424/B2 VGND VGND VPWR VPWR U$$1417/A sky130_fd_sc_hd__a22o_1
XFILLER_167_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1427 U$$1427/A U$$1459/B VGND VGND VPWR VPWR U$$1427/X sky130_fd_sc_hd__xor2_1
XU$$1438 U$$3354/B1 U$$1442/A2 U$$344/A1 U$$1442/B2 VGND VGND VPWR VPWR U$$1439/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1449 U$$1449/A U$$1487/B VGND VGND VPWR VPWR U$$1449/X sky130_fd_sc_hd__xor2_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_308 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_216_ _351_/CLK _216_/D VGND VGND VPWR VPWR _216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4253_1766 VGND VGND VPWR VPWR U$$4253_1766/HI U$$4253/A1 sky130_fd_sc_hd__conb_1
XFILLER_66_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_52_4 dadda_fa_2_52_4/A dadda_fa_2_52_4/B dadda_fa_2_52_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/CIN dadda_fa_3_52_3/CIN sky130_fd_sc_hd__fa_1
XU$$4020 U$$4020/A U$$4058/B VGND VGND VPWR VPWR U$$4020/X sky130_fd_sc_hd__xor2_1
XFILLER_39_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4031 U$$4442/A1 U$$4071/A2 U$$4031/B1 U$$4071/B2 VGND VGND VPWR VPWR U$$4032/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4042 U$$4042/A U$$4072/B VGND VGND VPWR VPWR U$$4042/X sky130_fd_sc_hd__xor2_1
XU$$4053 U$$4053/A1 U$$4061/A2 _589_/Q U$$4061/B2 VGND VGND VPWR VPWR U$$4054/A sky130_fd_sc_hd__a22o_1
XU$$4064 U$$4064/A U$$4070/B VGND VGND VPWR VPWR U$$4064/X sky130_fd_sc_hd__xor2_1
XFILLER_65_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_45_3 dadda_fa_2_45_3/A dadda_fa_2_45_3/B dadda_fa_2_45_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_1/B dadda_fa_3_45_3/B sky130_fd_sc_hd__fa_1
XU$$3330 U$$4426/A1 U$$3368/A2 _570_/Q U$$3368/B2 VGND VGND VPWR VPWR U$$3331/A sky130_fd_sc_hd__a22o_1
XU$$4075 U$$4075/A1 U$$3977/X U$$4351/A1 U$$3978/X VGND VGND VPWR VPWR U$$4076/A sky130_fd_sc_hd__a22o_1
XU$$4086 U$$4086/A U$$4109/A VGND VGND VPWR VPWR U$$4086/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3341 U$$3341/A U$$3343/B VGND VGND VPWR VPWR U$$3341/X sky130_fd_sc_hd__xor2_1
XU$$3352 U$$3352/A1 U$$3404/A2 U$$4450/A1 U$$3404/B2 VGND VGND VPWR VPWR U$$3353/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_38_2 U$$1945/X U$$2078/X U$$2211/X VGND VGND VPWR VPWR dadda_fa_3_39_1/A
+ dadda_fa_3_38_3/A sky130_fd_sc_hd__fa_1
XU$$4097 U$$4369/B1 U$$4107/A2 U$$4236/A1 U$$4105/B2 VGND VGND VPWR VPWR U$$4098/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3363 U$$3363/A U$$3363/B VGND VGND VPWR VPWR U$$3363/X sky130_fd_sc_hd__xor2_1
XU$$3374 U$$3374/A1 U$$3418/A2 U$$4472/A1 U$$3418/B2 VGND VGND VPWR VPWR U$$3375/A
+ sky130_fd_sc_hd__a22o_1
XU$$2640 U$$2640/A U$$2688/B VGND VGND VPWR VPWR U$$2640/X sky130_fd_sc_hd__xor2_1
XU$$3385 U$$3385/A U$$3397/B VGND VGND VPWR VPWR U$$3385/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_15_1 dadda_fa_5_15_1/A dadda_fa_5_15_1/B dadda_fa_5_15_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_16_0/B dadda_fa_7_15_0/A sky130_fd_sc_hd__fa_2
XU$$3396 U$$3805/B1 U$$3402/A2 _603_/Q U$$3402/B2 VGND VGND VPWR VPWR U$$3397/A sky130_fd_sc_hd__a22o_1
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2651 U$$2786/B1 U$$2653/A2 U$$3475/A1 U$$2653/B2 VGND VGND VPWR VPWR U$$2652/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2662 U$$2662/A U$$2664/B VGND VGND VPWR VPWR U$$2662/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2673 U$$3769/A1 U$$2707/A2 U$$3769/B1 U$$2707/B2 VGND VGND VPWR VPWR U$$2674/A
+ sky130_fd_sc_hd__a22o_1
XU$$2684 U$$2684/A U$$2688/B VGND VGND VPWR VPWR U$$2684/X sky130_fd_sc_hd__xor2_1
XFILLER_61_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2695 U$$3380/A1 U$$2733/A2 U$$368/A1 U$$2733/B2 VGND VGND VPWR VPWR U$$2696/A
+ sky130_fd_sc_hd__a22o_1
XU$$1950 U$$32/A1 U$$1956/A2 U$$34/A1 U$$1956/B2 VGND VGND VPWR VPWR U$$1951/A sky130_fd_sc_hd__a22o_1
XFILLER_210_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1961 U$$1961/A U$$2011/B VGND VGND VPWR VPWR U$$1961/X sky130_fd_sc_hd__xor2_1
XU$$1972 U$$3753/A1 U$$1976/A2 U$$3618/A1 U$$1976/B2 VGND VGND VPWR VPWR U$$1973/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1983 U$$1983/A U$$1983/B VGND VGND VPWR VPWR U$$1983/X sky130_fd_sc_hd__xor2_1
XU$$1994 U$$624/A1 U$$1922/X U$$624/B1 U$$1923/X VGND VGND VPWR VPWR U$$1995/A sky130_fd_sc_hd__a22o_1
XFILLER_166_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_371 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_859 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput108 b[49] VGND VGND VPWR VPWR _601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput119 b[59] VGND VGND VPWR VPWR _611_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$613 final_adder.U$$740/A final_adder.U$$740/B final_adder.U$$613/B1
+ VGND VGND VPWR VPWR final_adder.U$$741/B sky130_fd_sc_hd__a21o_1
XTAP_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$624 final_adder.U$$624/A final_adder.U$$624/B VGND VGND VPWR VPWR
+ _170_/D sky130_fd_sc_hd__xor2_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$635 final_adder.U$$635/A final_adder.U$$635/B VGND VGND VPWR VPWR
+ _181_/D sky130_fd_sc_hd__xor2_4
XFILLER_116_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater850 U$$1587/B2 VGND VGND VPWR VPWR U$$1577/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$646 final_adder.U$$646/A final_adder.U$$646/B VGND VGND VPWR VPWR
+ _192_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$657 final_adder.U$$657/A final_adder.U$$657/B VGND VGND VPWR VPWR
+ _203_/D sky130_fd_sc_hd__xor2_1
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater861 U$$259/B2 VGND VGND VPWR VPWR U$$217/B2 sky130_fd_sc_hd__buf_4
XFILLER_186_1003 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$507 U$$916/B1 U$$517/A2 U$$781/B1 U$$517/B2 VGND VGND VPWR VPWR U$$508/A sky130_fd_sc_hd__a22o_1
XFILLER_29_469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$668 final_adder.U$$668/A final_adder.U$$668/B VGND VGND VPWR VPWR
+ _214_/D sky130_fd_sc_hd__xor2_4
Xrepeater872 U$$1295/B2 VGND VGND VPWR VPWR U$$1279/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$679 final_adder.U$$679/A final_adder.U$$679/B VGND VGND VPWR VPWR
+ _225_/D sky130_fd_sc_hd__xor2_1
XU$$518 U$$518/A U$$518/B VGND VGND VPWR VPWR U$$518/X sky130_fd_sc_hd__xor2_1
Xrepeater883 U$$1194/B2 VGND VGND VPWR VPWR U$$1190/B2 sky130_fd_sc_hd__buf_4
XFILLER_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_40_2 U$$885/X U$$1018/X U$$1151/X VGND VGND VPWR VPWR dadda_fa_2_41_4/B
+ dadda_fa_2_40_5/CIN sky130_fd_sc_hd__fa_1
Xrepeater894 U$$5/X VGND VGND VPWR VPWR U$$98/B2 sky130_fd_sc_hd__buf_4
XU$$529 U$$938/B1 U$$415/X U$$805/A1 U$$416/X VGND VGND VPWR VPWR U$$530/A sky130_fd_sc_hd__a22o_1
XFILLER_38_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$90 U$$90/A1 U$$4/X U$$92/A1 U$$5/X VGND VGND VPWR VPWR U$$91/A sky130_fd_sc_hd__a22o_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_10_0 U$$27/X U$$160/X U$$293/X VGND VGND VPWR VPWR dadda_fa_5_11_0/CIN
+ dadda_fa_5_10_1/B sky130_fd_sc_hd__fa_1
XFILLER_188_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_70 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_81 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_92 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1407 _589_/Q VGND VGND VPWR VPWR U$$3916/B1 sky130_fd_sc_hd__buf_4
XFILLER_21_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1418 _588_/Q VGND VGND VPWR VPWR U$$4053/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_114_0 dadda_fa_3_114_0/A U$$3560/X U$$3693/X VGND VGND VPWR VPWR dadda_fa_4_115_2/A
+ dadda_fa_4_114_2/B sky130_fd_sc_hd__fa_1
XFILLER_119_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1429 U$$3362/B1 VGND VGND VPWR VPWR U$$896/B1 sky130_fd_sc_hd__buf_12
XFILLER_197_1187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_62_3 dadda_fa_3_62_3/A dadda_fa_3_62_3/B dadda_fa_3_62_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_1/B dadda_fa_4_62_2/CIN sky130_fd_sc_hd__fa_1
Xclkbuf_2_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_2_0_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_55_2 dadda_fa_3_55_2/A dadda_fa_3_55_2/B dadda_fa_3_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_1/A dadda_fa_4_55_2/B sky130_fd_sc_hd__fa_1
XFILLER_47_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_48_1 dadda_fa_3_48_1/A dadda_fa_3_48_1/B dadda_fa_3_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_0/CIN dadda_fa_4_48_2/A sky130_fd_sc_hd__fa_1
XFILLER_29_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_25_0 dadda_fa_6_25_0/A dadda_fa_6_25_0/B dadda_fa_6_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_26_0/B dadda_fa_7_25_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_90_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1202 U$$928/A1 U$$1100/X U$$930/A1 U$$1101/X VGND VGND VPWR VPWR U$$1203/A sky130_fd_sc_hd__a22o_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1213 U$$1213/A U$$1232/A VGND VGND VPWR VPWR U$$1213/X sky130_fd_sc_hd__xor2_1
XU$$1224 U$$948/B1 U$$1224/A2 U$$952/A1 U$$1224/B2 VGND VGND VPWR VPWR U$$1225/A sky130_fd_sc_hd__a22o_1
XU$$1235 U$$1370/A VGND VGND VPWR VPWR U$$1235/Y sky130_fd_sc_hd__inv_1
XFILLER_16_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1246 U$$1246/A U$$1280/B VGND VGND VPWR VPWR U$$1246/X sky130_fd_sc_hd__xor2_1
XFILLER_16_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1257 U$$435/A1 U$$1323/A2 U$$435/B1 U$$1323/B2 VGND VGND VPWR VPWR U$$1258/A sky130_fd_sc_hd__a22o_1
XFILLER_71_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1268 U$$1268/A U$$1280/B VGND VGND VPWR VPWR U$$1268/X sky130_fd_sc_hd__xor2_1
XFILLER_15_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1279 U$$46/A1 U$$1279/A2 U$$48/A1 U$$1279/B2 VGND VGND VPWR VPWR U$$1280/A sky130_fd_sc_hd__a22o_1
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_896 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_50_1 dadda_fa_2_50_1/A dadda_fa_2_50_1/B dadda_fa_2_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_0/CIN dadda_fa_3_50_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_22_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4411_1784 VGND VGND VPWR VPWR U$$4411_1784/HI U$$4411/B sky130_fd_sc_hd__conb_1
XFILLER_22_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_43_0 U$$1955/X U$$2088/X U$$2221/X VGND VGND VPWR VPWR dadda_fa_3_44_0/B
+ dadda_fa_3_43_2/B sky130_fd_sc_hd__fa_1
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3160 U$$3160/A U$$3208/B VGND VGND VPWR VPWR U$$3160/X sky130_fd_sc_hd__xor2_1
XU$$3171 U$$3445/A1 U$$3215/A2 U$$3310/A1 U$$3215/B2 VGND VGND VPWR VPWR U$$3172/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3182 U$$3182/A U$$3208/B VGND VGND VPWR VPWR U$$3182/X sky130_fd_sc_hd__xor2_1
XU$$3193 U$$3193/A1 U$$3235/A2 U$$4291/A1 U$$3235/B2 VGND VGND VPWR VPWR U$$3194/A
+ sky130_fd_sc_hd__a22o_1
XU$$2470 U$$2468/Y _652_/Q U$$2466/A U$$2469/X U$$2466/Y VGND VGND VPWR VPWR U$$2470/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_62_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2481 U$$2481/A U$$2541/B VGND VGND VPWR VPWR U$$2481/X sky130_fd_sc_hd__xor2_1
XFILLER_50_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2492 U$$985/A1 U$$2516/A2 U$$987/A1 U$$2516/B2 VGND VGND VPWR VPWR U$$2493/A sky130_fd_sc_hd__a22o_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1780 U$$1780/A VGND VGND VPWR VPWR U$$1780/Y sky130_fd_sc_hd__inv_1
XU$$1791 U$$969/A1 U$$1859/A2 U$$971/A1 U$$1859/B2 VGND VGND VPWR VPWR U$$1792/A sky130_fd_sc_hd__a22o_1
XFILLER_50_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 b[32] VGND VGND VPWR VPWR _584_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_72_2 dadda_fa_4_72_2/A dadda_fa_4_72_2/B dadda_fa_4_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/CIN dadda_fa_5_72_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_88_2 U$$2444/X U$$2577/X U$$2710/X VGND VGND VPWR VPWR dadda_fa_2_89_4/A
+ dadda_fa_2_88_5/B sky130_fd_sc_hd__fa_1
XFILLER_116_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_65_1 dadda_fa_4_65_1/A dadda_fa_4_65_1/B dadda_fa_4_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/B dadda_fa_5_65_1/B sky130_fd_sc_hd__fa_1
XFILLER_115_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_42_0 dadda_fa_7_42_0/A dadda_fa_7_42_0/B dadda_fa_7_42_0/CIN VGND VGND
+ VPWR VPWR _467_/D _338_/D sky130_fd_sc_hd__fa_1
XFILLER_103_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_58_0 dadda_fa_4_58_0/A dadda_fa_4_58_0/B dadda_fa_4_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/A dadda_fa_5_58_1/A sky130_fd_sc_hd__fa_1
XFILLER_88_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$421 final_adder.U$$338/B final_adder.U$$694/B final_adder.U$$293/X
+ VGND VGND VPWR VPWR final_adder.U$$698/B sky130_fd_sc_hd__a21o_1
XTAP_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$443 final_adder.U$$266/B final_adder.U$$642/B final_adder.U$$149/X
+ VGND VGND VPWR VPWR final_adder.U$$644/B sky130_fd_sc_hd__a21o_1
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$304 U$$30/A1 U$$334/A2 U$$991/A1 U$$334/B2 VGND VGND VPWR VPWR U$$305/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$465 final_adder.U$$288/B final_adder.U$$686/B final_adder.U$$193/X
+ VGND VGND VPWR VPWR final_adder.U$$688/B sky130_fd_sc_hd__a21o_1
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$315 U$$315/A U$$319/B VGND VGND VPWR VPWR U$$315/X sky130_fd_sc_hd__xor2_1
X_550_ _550_/CLK _550_/D VGND VGND VPWR VPWR _550_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater680 U$$457/B2 VGND VGND VPWR VPWR U$$447/B2 sky130_fd_sc_hd__buf_4
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$326 U$$463/A1 U$$334/A2 U$$463/B1 U$$334/B2 VGND VGND VPWR VPWR U$$327/A sky130_fd_sc_hd__a22o_1
XFILLER_72_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$487 final_adder.U$$310/B final_adder.U$$730/B final_adder.U$$237/X
+ VGND VGND VPWR VPWR final_adder.U$$732/B sky130_fd_sc_hd__a21o_1
Xrepeater691 U$$4115/X VGND VGND VPWR VPWR U$$4174/B2 sky130_fd_sc_hd__buf_6
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$337 U$$337/A U$$351/B VGND VGND VPWR VPWR U$$337/X sky130_fd_sc_hd__xor2_1
XFILLER_205_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_25 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$348 U$$896/A1 U$$350/A2 U$$898/A1 U$$350/B2 VGND VGND VPWR VPWR U$$349/A sky130_fd_sc_hd__a22o_1
XU$$359 U$$359/A U$$397/B VGND VGND VPWR VPWR U$$359/X sky130_fd_sc_hd__xor2_1
X_481_ _482_/CLK _481_/D VGND VGND VPWR VPWR _481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1204 U$$2459/B1 VGND VGND VPWR VPWR U$$954/A1 sky130_fd_sc_hd__buf_6
Xrepeater1215 _613_/Q VGND VGND VPWR VPWR U$$2459/A1 sky130_fd_sc_hd__buf_4
XFILLER_165_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1226 U$$946/B1 VGND VGND VPWR VPWR U$$811/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_5_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1237 U$$3412/A1 VGND VGND VPWR VPWR U$$4508/A1 sky130_fd_sc_hd__buf_4
XFILLER_114_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1248 U$$2721/B1 VGND VGND VPWR VPWR U$$942/A1 sky130_fd_sc_hd__clkbuf_8
Xrepeater1259 U$$4502/A1 VGND VGND VPWR VPWR U$$4500/B1 sky130_fd_sc_hd__buf_4
XFILLER_113_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_60_0 dadda_fa_3_60_0/A dadda_fa_3_60_0/B dadda_fa_3_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_0/B dadda_fa_4_60_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_76_0 dadda_fa_0_76_0/A U$$957/X U$$1090/X VGND VGND VPWR VPWR dadda_fa_1_77_8/B
+ dadda_fa_1_76_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$860 U$$38/A1 U$$860/A2 U$$40/A1 U$$860/B2 VGND VGND VPWR VPWR U$$861/A sky130_fd_sc_hd__a22o_1
XU$$1010 U$$1010/A U$$980/B VGND VGND VPWR VPWR U$$1010/X sky130_fd_sc_hd__xor2_1
XU$$871 U$$871/A U$$879/B VGND VGND VPWR VPWR U$$871/X sky130_fd_sc_hd__xor2_1
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_679_ _679_/CLK _679_/D VGND VGND VPWR VPWR _679_/Q sky130_fd_sc_hd__dfxtp_4
XU$$1021 U$$62/A1 U$$1065/A2 U$$64/A1 U$$1065/B2 VGND VGND VPWR VPWR U$$1022/A sky130_fd_sc_hd__a22o_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$882 U$$882/A1 U$$906/A2 U$$882/B1 U$$906/B2 VGND VGND VPWR VPWR U$$883/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$893 U$$893/A U$$925/B VGND VGND VPWR VPWR U$$893/X sky130_fd_sc_hd__xor2_1
XU$$1032 U$$1032/A U$$1040/B VGND VGND VPWR VPWR U$$1032/X sky130_fd_sc_hd__xor2_1
XFILLER_189_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1043 U$$906/A1 U$$1089/A2 U$$908/A1 U$$1089/B2 VGND VGND VPWR VPWR U$$1044/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1054 U$$1054/A U$$998/B VGND VGND VPWR VPWR U$$1054/X sky130_fd_sc_hd__xor2_1
XU$$1065 U$$928/A1 U$$1065/A2 U$$930/A1 U$$1065/B2 VGND VGND VPWR VPWR U$$1066/A sky130_fd_sc_hd__a22o_1
XFILLER_149_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1076 U$$1076/A U$$1078/B VGND VGND VPWR VPWR U$$1076/X sky130_fd_sc_hd__xor2_1
XFILLER_204_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1087 U$$948/B1 U$$1089/A2 U$$952/A1 U$$1089/B2 VGND VGND VPWR VPWR U$$1088/A sky130_fd_sc_hd__a22o_1
XU$$1098 _633_/Q VGND VGND VPWR VPWR U$$1098/Y sky130_fd_sc_hd__inv_1
XFILLER_188_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4441_1799 VGND VGND VPWR VPWR U$$4441_1799/HI U$$4441/B sky130_fd_sc_hd__conb_1
XFILLER_191_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_694 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_82_1 dadda_fa_5_82_1/A dadda_fa_5_82_1/B dadda_fa_5_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_83_0/B dadda_fa_7_82_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_98_1 U$$2730/X U$$2863/X U$$2996/X VGND VGND VPWR VPWR dadda_fa_3_99_1/A
+ dadda_fa_3_98_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4517_1837 VGND VGND VPWR VPWR U$$4517_1837/HI U$$4517/B sky130_fd_sc_hd__conb_1
XFILLER_7_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_75_0 dadda_fa_5_75_0/A dadda_fa_5_75_0/B dadda_fa_5_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_76_0/A dadda_fa_6_75_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_98_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_74_8 dadda_fa_1_74_8/A dadda_fa_1_74_8/B dadda_fa_1_74_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_75_3/A dadda_fa_3_74_0/A sky130_fd_sc_hd__fa_2
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_67_7 dadda_fa_1_67_7/A dadda_fa_1_67_7/B dadda_fa_1_67_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_2/CIN dadda_fa_2_67_5/CIN sky130_fd_sc_hd__fa_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_832 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1042 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_93_0 U$$2054/Y U$$2188/X U$$2321/X VGND VGND VPWR VPWR dadda_fa_2_94_5/A
+ dadda_fa_2_93_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_155_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3907 U$$3907/A U$$3933/B VGND VGND VPWR VPWR U$$3907/X sky130_fd_sc_hd__xor2_1
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$240 final_adder.U$$735/A ANTENNA_9/DIODE VGND VGND VPWR VPWR final_adder.U$$312/B
+ sky130_fd_sc_hd__and2_1
XU$$3918 _589_/Q U$$3932/A2 U$$4468/A1 U$$3932/B2 VGND VGND VPWR VPWR U$$3919/A sky130_fd_sc_hd__a22o_1
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$251 final_adder.U$$745/A final_adder.U$$617/B1 final_adder.U$$251/B1
+ VGND VGND VPWR VPWR final_adder.U$$251/X sky130_fd_sc_hd__a21o_1
X_602_ _613_/CLK _602_/D VGND VGND VPWR VPWR _602_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3929 U$$3929/A U$$3935/B VGND VGND VPWR VPWR U$$3929/X sky130_fd_sc_hd__xor2_1
XFILLER_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$101 U$$101/A U$$99/B VGND VGND VPWR VPWR U$$101/X sky130_fd_sc_hd__xor2_1
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$262 final_adder.U$$262/A final_adder.U$$262/B VGND VGND VPWR VPWR
+ final_adder.U$$322/A sky130_fd_sc_hd__and2_1
Xdadda_fa_6_105_0 dadda_fa_6_105_0/A dadda_fa_6_105_0/B dadda_fa_6_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_106_0/B dadda_fa_7_105_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$273 final_adder.U$$272/A final_adder.U$$161/X final_adder.U$$163/X
+ VGND VGND VPWR VPWR final_adder.U$$273/X sky130_fd_sc_hd__a21o_1
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$112 U$$384/B1 U$$118/A2 U$$251/A1 U$$118/B2 VGND VGND VPWR VPWR U$$113/A sky130_fd_sc_hd__a22o_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$284 final_adder.U$$284/A final_adder.U$$284/B VGND VGND VPWR VPWR
+ final_adder.U$$334/B sky130_fd_sc_hd__and2_1
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$123 U$$123/A U$$129/B VGND VGND VPWR VPWR U$$123/X sky130_fd_sc_hd__xor2_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$295 final_adder.U$$294/A final_adder.U$$205/X final_adder.U$$207/X
+ VGND VGND VPWR VPWR final_adder.U$$295/X sky130_fd_sc_hd__a21o_1
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$134 U$$406/B1 U$$4/X U$$134/B1 U$$5/X VGND VGND VPWR VPWR U$$135/A sky130_fd_sc_hd__a22o_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$145 U$$8/A1 U$$181/A2 U$$8/B1 U$$181/B2 VGND VGND VPWR VPWR U$$146/A sky130_fd_sc_hd__a22o_1
XFILLER_150_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_533_ _559_/CLK _533_/D VGND VGND VPWR VPWR _533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_25_3 dadda_fa_3_25_3/A dadda_fa_3_25_3/B dadda_fa_3_25_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_26_1/B dadda_fa_4_25_2/CIN sky130_fd_sc_hd__fa_1
XU$$156 U$$156/A U$$190/B VGND VGND VPWR VPWR U$$156/X sky130_fd_sc_hd__xor2_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$167 U$$989/A1 U$$195/A2 U$$991/A1 U$$195/B2 VGND VGND VPWR VPWR U$$168/A sky130_fd_sc_hd__a22o_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$178 U$$178/A U$$180/B VGND VGND VPWR VPWR U$$178/X sky130_fd_sc_hd__xor2_1
XFILLER_207_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$189 U$$600/A1 U$$219/A2 U$$54/A1 U$$219/B2 VGND VGND VPWR VPWR U$$190/A sky130_fd_sc_hd__a22o_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_464_ _466_/CLK _464_/D VGND VGND VPWR VPWR _464_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_395_ _526_/CLK _395_/D VGND VGND VPWR VPWR _395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_92_0 dadda_fa_6_92_0/A dadda_fa_6_92_0/B dadda_fa_6_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_93_0/B dadda_fa_7_92_0/CIN sky130_fd_sc_hd__fa_2
Xrepeater1001 U$$3014/A VGND VGND VPWR VPWR U$$2972/B sky130_fd_sc_hd__buf_6
XFILLER_86_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1012 U$$2708/B VGND VGND VPWR VPWR U$$2698/B sky130_fd_sc_hd__buf_8
Xrepeater1023 U$$2567/B VGND VGND VPWR VPWR U$$2541/B sky130_fd_sc_hd__buf_12
Xrepeater1034 U$$2400/B VGND VGND VPWR VPWR U$$2388/B sky130_fd_sc_hd__buf_6
XFILLER_86_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1045 U$$2309/B VGND VGND VPWR VPWR U$$2321/B sky130_fd_sc_hd__buf_6
Xrepeater1056 U$$2043/B VGND VGND VPWR VPWR U$$1957/B sky130_fd_sc_hd__buf_8
XFILLER_5_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1067 U$$1852/B VGND VGND VPWR VPWR U$$1844/B sky130_fd_sc_hd__buf_8
Xrepeater1078 U$$1747/B VGND VGND VPWR VPWR U$$1723/B sky130_fd_sc_hd__buf_12
Xrepeater1089 U$$1636/B VGND VGND VPWR VPWR U$$1628/B sky130_fd_sc_hd__buf_6
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$690 U$$688/B _625_/Q _626_/Q U$$685/Y VGND VGND VPWR VPWR U$$690/X sky130_fd_sc_hd__a22o_2
XFILLER_211_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_2__f_clk clkbuf_2_1_0_clk/X VGND VGND VPWR VPWR _432_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_80_8 U$$4290/X U$$4423/X VGND VGND VPWR VPWR dadda_fa_2_81_3/B dadda_fa_3_80_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1590 U$$310/A1 VGND VGND VPWR VPWR U$$719/B1 sky130_fd_sc_hd__buf_8
XFILLER_28_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_72_5 U$$4008/X U$$4141/X U$$4274/X VGND VGND VPWR VPWR dadda_fa_2_73_2/A
+ dadda_fa_2_72_5/A sky130_fd_sc_hd__fa_1
XFILLER_150_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_65_4 U$$4127/X U$$4260/X U$$4393/X VGND VGND VPWR VPWR dadda_fa_2_66_1/CIN
+ dadda_fa_2_65_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_82_0_1855 VGND VGND VPWR VPWR dadda_fa_1_82_0/A dadda_fa_1_82_0_1855/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_46_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_58_3 U$$2783/X U$$2916/X U$$3049/X VGND VGND VPWR VPWR dadda_fa_2_59_1/B
+ dadda_fa_2_58_4/B sky130_fd_sc_hd__fa_1
XFILLER_100_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_35_2 dadda_fa_4_35_2/A dadda_fa_4_35_2/B dadda_fa_4_35_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/CIN dadda_fa_5_35_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_28_1 dadda_fa_4_28_1/A dadda_fa_4_28_1/B dadda_fa_4_28_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/B dadda_fa_5_28_1/B sky130_fd_sc_hd__fa_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_180_ _189_/CLK _180_/D VGND VGND VPWR VPWR _180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_79 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4405 U$$4405/A U$$4405/B VGND VGND VPWR VPWR U$$4405/X sky130_fd_sc_hd__xor2_1
XU$$4416 U$$4416/A1 U$$4388/X U$$4418/A1 U$$4430/B2 VGND VGND VPWR VPWR U$$4417/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_60_3 U$$1324/X U$$1457/X U$$1590/X VGND VGND VPWR VPWR dadda_fa_1_61_7/A
+ dadda_fa_1_60_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4427 U$$4427/A U$$4427/B VGND VGND VPWR VPWR U$$4427/X sky130_fd_sc_hd__xor2_1
XFILLER_65_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4438 _575_/Q U$$4388/X U$$4440/A1 U$$4438/B2 VGND VGND VPWR VPWR U$$4439/A sky130_fd_sc_hd__a22o_1
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4449 U$$4449/A U$$4449/B VGND VGND VPWR VPWR U$$4449/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_17_1 U$$440/X U$$573/X VGND VGND VPWR VPWR dadda_fa_4_18_1/CIN dadda_ha_3_17_1/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_38_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3704 U$$3702/B U$$3699/A _670_/Q U$$3699/Y VGND VGND VPWR VPWR U$$3704/X sky130_fd_sc_hd__a22o_4
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3715 U$$4400/A1 U$$3769/A2 _557_/Q U$$3769/B2 VGND VGND VPWR VPWR U$$3716/A sky130_fd_sc_hd__a22o_1
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3726 U$$3726/A U$$3832/B VGND VGND VPWR VPWR U$$3726/X sky130_fd_sc_hd__xor2_1
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3737 U$$584/B1 U$$3743/A2 U$$451/A1 U$$3743/B2 VGND VGND VPWR VPWR U$$3738/A sky130_fd_sc_hd__a22o_1
XU$$3748 U$$3748/A U$$3760/B VGND VGND VPWR VPWR U$$3748/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_30_1 input180/X dadda_fa_3_30_1/B dadda_fa_3_30_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_31_0/CIN dadda_fa_4_30_2/A sky130_fd_sc_hd__fa_2
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3759 U$$4031/B1 U$$3777/A2 U$$3896/B1 U$$3777/B2 VGND VGND VPWR VPWR U$$3760/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1023 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_330 _239_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_23_0 U$$319/X U$$452/X U$$585/X VGND VGND VPWR VPWR dadda_fa_4_24_0/B
+ dadda_fa_4_23_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_341 U$$229/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_516_ _516_/CLK _516_/D VGND VGND VPWR VPWR _516_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_352 _638_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_363 _623_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_374 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_385 _648_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_447_ _448_/CLK _447_/D VGND VGND VPWR VPWR _447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_378_ _516_/CLK _378_/D VGND VGND VPWR VPWR _378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_336 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_82_4 dadda_fa_2_82_4/A dadda_fa_2_82_4/B dadda_fa_2_82_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/CIN dadda_fa_3_82_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_173_1027 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_75_3 dadda_fa_2_75_3/A dadda_fa_2_75_3/B dadda_fa_2_75_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/B dadda_fa_3_75_3/B sky130_fd_sc_hd__fa_1
XFILLER_141_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_68_2 dadda_fa_2_68_2/A dadda_fa_2_68_2/B dadda_fa_2_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/A dadda_fa_3_68_3/A sky130_fd_sc_hd__fa_2
XFILLER_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_70_0_1850 VGND VGND VPWR VPWR dadda_fa_0_70_0/A dadda_fa_0_70_0_1850/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_84_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_45_1 dadda_fa_5_45_1/A dadda_fa_5_45_1/B dadda_fa_5_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_46_0/B dadda_fa_7_45_0/A sky130_fd_sc_hd__fa_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_810 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_38_0 dadda_fa_5_38_0/A dadda_fa_5_38_0/B dadda_fa_5_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_39_0/A dadda_fa_6_38_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_52_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_112_0 dadda_fa_5_112_0/A dadda_fa_5_112_0/B dadda_fa_5_112_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_113_0/A dadda_fa_6_112_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_70_2 U$$3073/X U$$3206/X U$$3339/X VGND VGND VPWR VPWR dadda_fa_2_71_1/A
+ dadda_fa_2_70_4/A sky130_fd_sc_hd__fa_1
XFILLER_120_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_1 U$$2793/X U$$2926/X U$$3059/X VGND VGND VPWR VPWR dadda_fa_2_64_0/CIN
+ dadda_fa_2_63_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_40_0 dadda_fa_4_40_0/A dadda_fa_4_40_0/B dadda_fa_4_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/A dadda_fa_5_40_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_56_0 U$$1183/X U$$1316/X U$$1449/X VGND VGND VPWR VPWR dadda_fa_2_57_0/B
+ dadda_fa_2_56_3/B sky130_fd_sc_hd__fa_1
XFILLER_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1609 U$$924/A1 U$$1635/A2 U$$924/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1610/A sky130_fd_sc_hd__a22o_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_301_ _431_/CLK _301_/D VGND VGND VPWR VPWR _301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_232_ _234_/CLK _232_/D VGND VGND VPWR VPWR _232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_275 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_92_3 dadda_fa_3_92_3/A dadda_fa_3_92_3/B dadda_fa_3_92_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_1/B dadda_fa_4_92_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_85_2 dadda_fa_3_85_2/A dadda_fa_3_85_2/B dadda_fa_3_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_1/A dadda_fa_4_85_2/B sky130_fd_sc_hd__fa_1
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_78_1 dadda_fa_3_78_1/A dadda_fa_3_78_1/B dadda_fa_3_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_0/CIN dadda_fa_4_78_2/A sky130_fd_sc_hd__fa_1
XFILLER_123_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_55_0 dadda_fa_6_55_0/A dadda_fa_6_55_0/B dadda_fa_6_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_56_0/B dadda_fa_7_55_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater509 U$$3148/A2 VGND VGND VPWR VPWR U$$3144/A2 sky130_fd_sc_hd__buf_4
XU$$4202 U$$4337/B1 U$$4202/A2 _595_/Q U$$4202/B2 VGND VGND VPWR VPWR U$$4203/A sky130_fd_sc_hd__a22o_1
XU$$4213 U$$4213/A U$$4247/A VGND VGND VPWR VPWR U$$4213/X sky130_fd_sc_hd__xor2_1
XU$$4224 U$$4224/A1 U$$4226/A2 U$$4361/B1 U$$4226/B2 VGND VGND VPWR VPWR U$$4225/A
+ sky130_fd_sc_hd__a22o_1
XU$$4235 U$$4235/A U$$4239/B VGND VGND VPWR VPWR U$$4235/X sky130_fd_sc_hd__xor2_1
XU$$3501 U$$3638/A1 U$$3545/A2 U$$3503/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3502/A
+ sky130_fd_sc_hd__a22o_1
XU$$4246 U$$4246/A VGND VGND VPWR VPWR U$$4246/Y sky130_fd_sc_hd__inv_1
XFILLER_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4257 U$$4394/A1 U$$4297/A2 U$$4396/A1 U$$4297/B2 VGND VGND VPWR VPWR U$$4258/A
+ sky130_fd_sc_hd__a22o_1
XU$$3512 U$$3512/A U$$3562/A VGND VGND VPWR VPWR U$$3512/X sky130_fd_sc_hd__xor2_1
XU$$3523 _597_/Q U$$3531/A2 _598_/Q U$$3531/B2 VGND VGND VPWR VPWR U$$3524/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_114_2 dadda_fa_4_114_2/A dadda_fa_4_114_2/B dadda_ha_3_114_1/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_115_0/CIN dadda_fa_5_114_1/CIN sky130_fd_sc_hd__fa_1
XU$$4268 U$$4268/A U$$4298/B VGND VGND VPWR VPWR U$$4268/X sky130_fd_sc_hd__xor2_1
XU$$4279 U$$4416/A1 U$$4311/A2 U$$4418/A1 U$$4319/B2 VGND VGND VPWR VPWR U$$4280/A
+ sky130_fd_sc_hd__a22o_1
XU$$3534 U$$3534/A U$$3538/B VGND VGND VPWR VPWR U$$3534/X sky130_fd_sc_hd__xor2_1
XFILLER_46_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2800 U$$4168/B1 U$$2744/X U$$4035/A1 U$$2745/X VGND VGND VPWR VPWR U$$2801/A sky130_fd_sc_hd__a22o_1
XU$$3545 U$$4228/B1 U$$3545/A2 U$$4369/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3546/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2811 U$$2811/A U$$2813/B VGND VGND VPWR VPWR U$$2811/X sky130_fd_sc_hd__xor2_1
XU$$3556 U$$3556/A U$$3556/B VGND VGND VPWR VPWR U$$3556/X sky130_fd_sc_hd__xor2_1
XFILLER_34_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_107_1 dadda_fa_4_107_1/A dadda_fa_4_107_1/B dadda_fa_4_107_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/B dadda_fa_5_107_1/B sky130_fd_sc_hd__fa_1
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2822 U$$3916/B1 U$$2856/A2 U$$3783/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2823/A
+ sky130_fd_sc_hd__a22o_1
XU$$3567 U$$3565/B U$$3562/A _668_/Q U$$3562/Y VGND VGND VPWR VPWR U$$3567/X sky130_fd_sc_hd__a22o_2
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2833 U$$2833/A U$$2843/B VGND VGND VPWR VPWR U$$2833/X sky130_fd_sc_hd__xor2_1
XU$$3578 U$$3578/A1 U$$3612/A2 U$$3578/B1 U$$3612/B2 VGND VGND VPWR VPWR U$$3579/A
+ sky130_fd_sc_hd__a22o_1
XU$$3589 U$$3589/A U$$3609/B VGND VGND VPWR VPWR U$$3589/X sky130_fd_sc_hd__xor2_1
XU$$2844 U$$3529/A1 U$$2874/A2 U$$3942/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2845/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2855 U$$2855/A U$$2861/B VGND VGND VPWR VPWR U$$2855/X sky130_fd_sc_hd__xor2_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2866 U$$2866/A1 U$$2866/A2 U$$3005/A1 U$$2866/B2 VGND VGND VPWR VPWR U$$2867/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2877 U$$2877/A VGND VGND VPWR VPWR U$$2877/Y sky130_fd_sc_hd__inv_1
XANTENNA_160 _180_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2888 U$$2888/A U$$2928/B VGND VGND VPWR VPWR U$$2888/X sky130_fd_sc_hd__xor2_1
XU$$2899 U$$3310/A1 U$$2915/A2 U$$3175/A1 U$$2915/B2 VGND VGND VPWR VPWR U$$2900/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_182 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_193 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_80_1 dadda_fa_2_80_1/A dadda_fa_2_80_1/B dadda_fa_2_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_0/CIN dadda_fa_3_80_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_73_0 dadda_fa_2_73_0/A dadda_fa_2_73_0/B dadda_fa_2_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_0/B dadda_fa_3_73_2/B sky130_fd_sc_hd__fa_1
XFILLER_170_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_95_1 dadda_fa_4_95_1/A dadda_fa_4_95_1/B dadda_fa_4_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/B dadda_fa_5_95_1/B sky130_fd_sc_hd__fa_1
XFILLER_118_450 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_72_0 dadda_fa_7_72_0/A dadda_fa_7_72_0/B dadda_fa_7_72_0/CIN VGND VGND
+ VPWR VPWR _497_/D _368_/D sky130_fd_sc_hd__fa_1
XFILLER_152_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_88_0 dadda_fa_4_88_0/A dadda_fa_4_88_0/B dadda_fa_4_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/A dadda_fa_5_88_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_109_3 U$$4348/X U$$4481/X input139/X VGND VGND VPWR VPWR dadda_fa_4_110_1/B
+ dadda_fa_4_109_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_145_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput370 _255_/Q VGND VGND VPWR VPWR o[87] sky130_fd_sc_hd__buf_2
XFILLER_117_1028 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput381 _265_/Q VGND VGND VPWR VPWR o[97] sky130_fd_sc_hd__buf_2
XFILLER_156_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2107 U$$3751/A1 U$$2109/A2 U$$3753/A1 U$$2109/B2 VGND VGND VPWR VPWR U$$2108/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2118 U$$2118/A U$$2144/B VGND VGND VPWR VPWR U$$2118/X sky130_fd_sc_hd__xor2_1
XU$$2129 U$$759/A1 U$$2129/A2 U$$624/A1 U$$2129/B2 VGND VGND VPWR VPWR U$$2130/A sky130_fd_sc_hd__a22o_1
XFILLER_62_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_835 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1406 U$$2774/B1 U$$1442/A2 U$$2641/A1 U$$1442/B2 VGND VGND VPWR VPWR U$$1407/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1417 U$$1417/A U$$1425/B VGND VGND VPWR VPWR U$$1417/X sky130_fd_sc_hd__xor2_1
XU$$1428 U$$3346/A1 U$$1428/A2 U$$882/A1 U$$1428/B2 VGND VGND VPWR VPWR U$$1429/A
+ sky130_fd_sc_hd__a22o_1
XU$$1439 U$$1439/A U$$1443/B VGND VGND VPWR VPWR U$$1439/X sky130_fd_sc_hd__xor2_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_315 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_215_ _476_/CLK _215_/D VGND VGND VPWR VPWR _215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_90_0 dadda_fa_3_90_0/A dadda_fa_3_90_0/B dadda_fa_3_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_0/B dadda_fa_4_90_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_171_537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_52_5 dadda_fa_2_52_5/A dadda_fa_2_52_5/B dadda_fa_2_52_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_2/A dadda_fa_4_52_0/A sky130_fd_sc_hd__fa_1
XU$$4010 U$$4010/A U$$4044/B VGND VGND VPWR VPWR U$$4010/X sky130_fd_sc_hd__xor2_1
XU$$4021 U$$4156/B1 U$$4029/A2 U$$4160/A1 U$$4029/B2 VGND VGND VPWR VPWR U$$4022/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4032 U$$4032/A U$$4072/B VGND VGND VPWR VPWR U$$4032/X sky130_fd_sc_hd__xor2_1
XFILLER_38_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4043 U$$4180/A1 U$$4065/A2 U$$4045/A1 U$$4065/B2 VGND VGND VPWR VPWR U$$4044/A
+ sky130_fd_sc_hd__a22o_1
XU$$4054 U$$4054/A U$$4058/B VGND VGND VPWR VPWR U$$4054/X sky130_fd_sc_hd__xor2_1
XFILLER_76_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3320 U$$3320/A1 U$$3320/A2 U$$3320/B1 U$$3320/B2 VGND VGND VPWR VPWR U$$3321/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_45_4 dadda_fa_2_45_4/A dadda_fa_2_45_4/B dadda_fa_2_45_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_1/CIN dadda_fa_3_45_3/CIN sky130_fd_sc_hd__fa_1
XU$$4065 _594_/Q U$$4065/A2 U$$4065/B1 U$$4065/B2 VGND VGND VPWR VPWR U$$4066/A sky130_fd_sc_hd__a22o_1
XFILLER_47_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3331 U$$3331/A U$$3369/B VGND VGND VPWR VPWR U$$3331/X sky130_fd_sc_hd__xor2_1
XU$$4076 U$$4076/A U$$4084/B VGND VGND VPWR VPWR U$$4076/X sky130_fd_sc_hd__xor2_1
XU$$4087 U$$4087/A1 U$$4107/A2 U$$4087/B1 U$$4107/B2 VGND VGND VPWR VPWR U$$4088/A
+ sky130_fd_sc_hd__a22o_1
XU$$3342 U$$3342/A1 U$$3378/A2 U$$4027/B1 U$$3378/B2 VGND VGND VPWR VPWR U$$3343/A
+ sky130_fd_sc_hd__a22o_1
XU$$3353 U$$3353/A U$$3357/B VGND VGND VPWR VPWR U$$3353/X sky130_fd_sc_hd__xor2_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4098 U$$4098/A U$$4109/A VGND VGND VPWR VPWR U$$4098/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3364 U$$4323/A1 U$$3378/A2 U$$4462/A1 U$$3378/B2 VGND VGND VPWR VPWR U$$3365/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_38_3 U$$2344/X U$$2477/X U$$2610/X VGND VGND VPWR VPWR dadda_fa_3_39_1/B
+ dadda_fa_3_38_3/B sky130_fd_sc_hd__fa_1
XU$$2630 U$$2630/A U$$2698/B VGND VGND VPWR VPWR U$$2630/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3375 U$$3375/A U$$3407/B VGND VGND VPWR VPWR U$$3375/X sky130_fd_sc_hd__xor2_1
XFILLER_207_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2641 U$$2641/A1 U$$2687/A2 U$$2641/B1 U$$2687/B2 VGND VGND VPWR VPWR U$$2642/A
+ sky130_fd_sc_hd__a22o_1
XU$$3386 U$$3521/B1 U$$3404/A2 U$$3386/B1 U$$3404/B2 VGND VGND VPWR VPWR U$$3387/A
+ sky130_fd_sc_hd__a22o_1
XU$$3397 U$$3397/A U$$3397/B VGND VGND VPWR VPWR U$$3397/X sky130_fd_sc_hd__xor2_1
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2652 U$$2652/A U$$2654/B VGND VGND VPWR VPWR U$$2652/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2663 U$$4168/B1 U$$2663/A2 U$$4035/A1 U$$2663/B2 VGND VGND VPWR VPWR U$$2664/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2674 U$$2674/A U$$2708/B VGND VGND VPWR VPWR U$$2674/X sky130_fd_sc_hd__xor2_1
XU$$2685 U$$3916/B1 U$$2687/A2 U$$3783/A1 U$$2687/B2 VGND VGND VPWR VPWR U$$2686/A
+ sky130_fd_sc_hd__a22o_1
XU$$1940 U$$20/B1 U$$1976/A2 U$$2077/B1 U$$1976/B2 VGND VGND VPWR VPWR U$$1941/A sky130_fd_sc_hd__a22o_1
XU$$1951 U$$1951/A U$$1957/B VGND VGND VPWR VPWR U$$1951/X sky130_fd_sc_hd__xor2_1
XU$$2696 U$$2696/A U$$2734/B VGND VGND VPWR VPWR U$$2696/X sky130_fd_sc_hd__xor2_1
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1962 U$$44/A1 U$$2010/A2 U$$46/A1 U$$2010/B2 VGND VGND VPWR VPWR U$$1963/A sky130_fd_sc_hd__a22o_1
XU$$1973 U$$1973/A U$$1977/B VGND VGND VPWR VPWR U$$1973/X sky130_fd_sc_hd__xor2_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1984 U$$3626/B1 U$$2010/A2 U$$3493/A1 U$$2010/B2 VGND VGND VPWR VPWR U$$1985/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1995 U$$1995/A U$$2003/B VGND VGND VPWR VPWR U$$1995/X sky130_fd_sc_hd__xor2_1
XFILLER_147_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput109 b[4] VGND VGND VPWR VPWR _556_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$603 final_adder.U$$730/A final_adder.U$$730/B final_adder.U$$603/B1
+ VGND VGND VPWR VPWR final_adder.U$$731/B sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$625 final_adder.U$$625/A final_adder.U$$625/B VGND VGND VPWR VPWR
+ _171_/D sky130_fd_sc_hd__xor2_1
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$636 final_adder.U$$636/A final_adder.U$$636/B VGND VGND VPWR VPWR
+ _182_/D sky130_fd_sc_hd__xor2_4
Xrepeater840 U$$1649/X VGND VGND VPWR VPWR U$$1736/B2 sky130_fd_sc_hd__buf_4
XFILLER_96_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$647 final_adder.U$$647/A final_adder.U$$647/B VGND VGND VPWR VPWR
+ _193_/D sky130_fd_sc_hd__xor2_4
Xrepeater851 U$$1587/B2 VGND VGND VPWR VPWR U$$1561/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$658 final_adder.U$$658/A final_adder.U$$658/B VGND VGND VPWR VPWR
+ _204_/D sky130_fd_sc_hd__xor2_1
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater862 U$$263/B2 VGND VGND VPWR VPWR U$$259/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_186_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$508 U$$508/A U$$518/B VGND VGND VPWR VPWR U$$508/X sky130_fd_sc_hd__xor2_1
XFILLER_45_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$669 final_adder.U$$669/A final_adder.U$$669/B VGND VGND VPWR VPWR
+ _215_/D sky130_fd_sc_hd__xor2_4
Xrepeater873 U$$1295/B2 VGND VGND VPWR VPWR U$$1309/B2 sky130_fd_sc_hd__buf_4
Xrepeater884 U$$1208/B2 VGND VGND VPWR VPWR U$$1194/B2 sky130_fd_sc_hd__buf_4
XU$$519 U$$791/B1 U$$545/A2 U$$658/A1 U$$545/B2 VGND VGND VPWR VPWR U$$520/A sky130_fd_sc_hd__a22o_1
Xrepeater895 U$$5/X VGND VGND VPWR VPWR U$$62/B2 sky130_fd_sc_hd__buf_2
XFILLER_44_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$80 U$$80/A1 U$$84/A2 U$$80/B1 U$$84/B2 VGND VGND VPWR VPWR U$$81/A sky130_fd_sc_hd__a22o_1
XU$$91 U$$91/A U$$93/B VGND VGND VPWR VPWR U$$91/X sky130_fd_sc_hd__xor2_1
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1062 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_60 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_82 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_93 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1408 U$$3779/B1 VGND VGND VPWR VPWR U$$3505/B1 sky130_fd_sc_hd__buf_6
XFILLER_115_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1419 U$$3229/A1 VGND VGND VPWR VPWR U$$78/A1 sky130_fd_sc_hd__buf_4
XFILLER_107_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_107_0 U$$3413/X U$$3546/X U$$3679/X VGND VGND VPWR VPWR dadda_fa_4_108_0/B
+ dadda_fa_4_107_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_55_3 dadda_fa_3_55_3/A dadda_fa_3_55_3/B dadda_fa_3_55_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_1/B dadda_fa_4_55_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_48_2 dadda_fa_3_48_2/A dadda_fa_3_48_2/B dadda_fa_3_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_1/A dadda_fa_4_48_2/B sky130_fd_sc_hd__fa_1
XFILLER_78_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_18_0 dadda_fa_6_18_0/A dadda_fa_6_18_0/B dadda_fa_6_18_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_19_0/B dadda_fa_7_18_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1203 U$$1203/A U$$1203/B VGND VGND VPWR VPWR U$$1203/X sky130_fd_sc_hd__xor2_1
XU$$1214 U$$253/B1 U$$1224/A2 U$$942/A1 U$$1224/B2 VGND VGND VPWR VPWR U$$1215/A sky130_fd_sc_hd__a22o_1
XU$$1225 U$$1225/A U$$1225/B VGND VGND VPWR VPWR U$$1225/X sky130_fd_sc_hd__xor2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1236 U$$1370/A U$$1236/B VGND VGND VPWR VPWR U$$1236/X sky130_fd_sc_hd__and2_1
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1247 U$$2343/A1 U$$1295/A2 U$$16/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1248/A sky130_fd_sc_hd__a22o_1
XU$$1258 U$$1258/A U$$1288/B VGND VGND VPWR VPWR U$$1258/X sky130_fd_sc_hd__xor2_1
XFILLER_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1269 U$$2774/B1 U$$1279/A2 U$$2641/A1 U$$1279/B2 VGND VGND VPWR VPWR U$$1270/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_104_clk _616_/CLK VGND VGND VPWR VPWR _492_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_50_2 dadda_fa_2_50_2/A dadda_fa_2_50_2/B dadda_fa_2_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/A dadda_fa_3_50_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_43_1 U$$2354/X U$$2487/X U$$2620/X VGND VGND VPWR VPWR dadda_fa_3_44_0/CIN
+ dadda_fa_3_43_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_20_0 dadda_fa_5_20_0/A dadda_fa_5_20_0/B dadda_fa_5_20_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_21_0/A dadda_fa_6_20_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_36_0 U$$744/X U$$877/X U$$1010/X VGND VGND VPWR VPWR dadda_fa_3_37_0/B
+ dadda_fa_3_36_2/B sky130_fd_sc_hd__fa_1
XU$$3150 _661_/Q VGND VGND VPWR VPWR U$$3150/Y sky130_fd_sc_hd__inv_1
XFILLER_53_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3161 U$$3709/A1 U$$3209/A2 U$$3437/A1 U$$3209/B2 VGND VGND VPWR VPWR U$$3162/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_198_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3172 U$$3172/A U$$3218/B VGND VGND VPWR VPWR U$$3172/X sky130_fd_sc_hd__xor2_1
XU$$3183 U$$3320/A1 U$$3209/A2 U$$4007/A1 U$$3209/B2 VGND VGND VPWR VPWR U$$3184/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3194 U$$3194/A U$$3236/B VGND VGND VPWR VPWR U$$3194/X sky130_fd_sc_hd__xor2_1
XFILLER_179_412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2460 U$$2460/A U$$2462/B VGND VGND VPWR VPWR U$$2460/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2471 U$$2469/B _651_/Q _652_/Q U$$2466/Y VGND VGND VPWR VPWR U$$2471/X sky130_fd_sc_hd__a22o_4
XU$$2482 U$$2756/A1 U$$2530/A2 U$$2756/B1 U$$2530/B2 VGND VGND VPWR VPWR U$$2483/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2493 U$$2493/A U$$2541/B VGND VGND VPWR VPWR U$$2493/X sky130_fd_sc_hd__xor2_1
XFILLER_179_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1770 U$$811/A1 U$$1778/A2 U$$950/A1 U$$1778/B2 VGND VGND VPWR VPWR U$$1771/A sky130_fd_sc_hd__a22o_1
XFILLER_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1781 _641_/Q VGND VGND VPWR VPWR U$$1781/Y sky130_fd_sc_hd__inv_1
XFILLER_72_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1792 U$$1792/A U$$1820/B VGND VGND VPWR VPWR U$$1792/X sky130_fd_sc_hd__xor2_1
XFILLER_50_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput80 b[23] VGND VGND VPWR VPWR _575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput91 b[33] VGND VGND VPWR VPWR _585_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_88_3 U$$2843/X U$$2976/X U$$3109/X VGND VGND VPWR VPWR dadda_fa_2_89_4/B
+ dadda_fa_2_88_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_153_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_65_2 dadda_fa_4_65_2/A dadda_fa_4_65_2/B dadda_fa_4_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/CIN dadda_fa_5_65_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_58_1 dadda_fa_4_58_1/A dadda_fa_4_58_1/B dadda_fa_4_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/B dadda_fa_5_58_1/B sky130_fd_sc_hd__fa_1
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$411 final_adder.U$$328/B final_adder.U$$654/B final_adder.U$$273/X
+ VGND VGND VPWR VPWR final_adder.U$$658/B sky130_fd_sc_hd__a21o_1
Xdadda_fa_7_35_0 dadda_fa_7_35_0/A dadda_fa_7_35_0/B dadda_fa_7_35_0/CIN VGND VGND
+ VPWR VPWR _460_/D _331_/D sky130_fd_sc_hd__fa_1
XTAP_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$433 final_adder.U$$316/X final_adder.U$$742/B final_adder.U$$317/X
+ VGND VGND VPWR VPWR final_adder.U$$746/B sky130_fd_sc_hd__a21o_2
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$455 final_adder.U$$278/B final_adder.U$$666/B final_adder.U$$173/X
+ VGND VGND VPWR VPWR final_adder.U$$668/B sky130_fd_sc_hd__a21o_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$305 U$$305/A U$$335/B VGND VGND VPWR VPWR U$$305/X sky130_fd_sc_hd__xor2_1
Xrepeater670 U$$553/X VGND VGND VPWR VPWR U$$682/B2 sky130_fd_sc_hd__buf_6
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater681 U$$491/B2 VGND VGND VPWR VPWR U$$457/B2 sky130_fd_sc_hd__clkbuf_4
Xfinal_adder.U$$477 final_adder.U$$300/B final_adder.U$$710/B final_adder.U$$217/X
+ VGND VGND VPWR VPWR final_adder.U$$712/B sky130_fd_sc_hd__a21o_1
XU$$316 U$$316/A1 U$$350/A2 U$$44/A1 U$$350/B2 VGND VGND VPWR VPWR U$$317/A sky130_fd_sc_hd__a22o_1
Xrepeater692 U$$4196/B2 VGND VGND VPWR VPWR U$$4182/B2 sky130_fd_sc_hd__buf_4
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$327 U$$327/A U$$335/B VGND VGND VPWR VPWR U$$327/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$499 final_adder.U$$626/A final_adder.U$$626/B final_adder.U$$499/B1
+ VGND VGND VPWR VPWR final_adder.U$$627/B sky130_fd_sc_hd__a21o_1
XU$$338 U$$747/B1 U$$350/A2 U$$614/A1 U$$350/B2 VGND VGND VPWR VPWR U$$339/A sky130_fd_sc_hd__a22o_1
XFILLER_38_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$349 U$$349/A U$$351/B VGND VGND VPWR VPWR U$$349/X sky130_fd_sc_hd__xor2_1
X_480_ _482_/CLK _480_/D VGND VGND VPWR VPWR _480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4427_1792 VGND VGND VPWR VPWR U$$4427_1792/HI U$$4427/B sky130_fd_sc_hd__conb_1
XFILLER_158_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1205 U$$3283/A1 VGND VGND VPWR VPWR U$$4516/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_148_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1216 U$$950/A1 VGND VGND VPWR VPWR U$$676/A1 sky130_fd_sc_hd__buf_4
XFILLER_181_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1227 U$$2866/A1 VGND VGND VPWR VPWR U$$946/B1 sky130_fd_sc_hd__buf_6
Xrepeater1238 U$$2999/B1 VGND VGND VPWR VPWR U$$3412/A1 sky130_fd_sc_hd__buf_6
Xrepeater1249 _608_/Q VGND VGND VPWR VPWR U$$2721/B1 sky130_fd_sc_hd__buf_6
XFILLER_84_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_60_1 dadda_fa_3_60_1/A dadda_fa_3_60_1/B dadda_fa_3_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_0/CIN dadda_fa_4_60_2/A sky130_fd_sc_hd__fa_1
XFILLER_122_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_53_0 dadda_fa_3_53_0/A dadda_fa_3_53_0/B dadda_fa_3_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_0/B dadda_fa_4_53_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_209_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_69_0 U$$410/Y U$$544/X U$$677/X VGND VGND VPWR VPWR dadda_fa_1_70_6/A
+ dadda_fa_1_69_7/CIN sky130_fd_sc_hd__fa_1
XU$$828_1845 VGND VGND VPWR VPWR U$$828_1845/HI U$$828/A1 sky130_fd_sc_hd__conb_1
XTAP_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$850 U$$28/A1 U$$924/A2 U$$30/A1 U$$924/B2 VGND VGND VPWR VPWR U$$851/A sky130_fd_sc_hd__a22o_1
X_678_ _679_/CLK _678_/D VGND VGND VPWR VPWR _678_/Q sky130_fd_sc_hd__dfxtp_1
XU$$861 U$$861/A U$$929/B VGND VGND VPWR VPWR U$$861/X sky130_fd_sc_hd__xor2_1
XU$$1000 U$$999/X U$$982/B VGND VGND VPWR VPWR U$$1000/X sky130_fd_sc_hd__xor2_1
XU$$872 U$$48/B1 U$$878/A2 U$$874/A1 U$$878/B2 VGND VGND VPWR VPWR U$$873/A sky130_fd_sc_hd__a22o_1
XU$$1011 U$$874/A1 U$$979/A2 U$$876/A1 U$$979/B2 VGND VGND VPWR VPWR U$$1012/A sky130_fd_sc_hd__a22o_1
XU$$1022 U$$1022/A U$$996/B VGND VGND VPWR VPWR U$$1022/X sky130_fd_sc_hd__xor2_1
XU$$883 U$$883/A U$$907/B VGND VGND VPWR VPWR U$$883/X sky130_fd_sc_hd__xor2_1
XU$$894 U$$894/A1 U$$896/A2 U$$896/A1 U$$896/B2 VGND VGND VPWR VPWR U$$895/A sky130_fd_sc_hd__a22o_1
XU$$1033 U$$896/A1 U$$1039/A2 U$$898/A1 U$$1039/B2 VGND VGND VPWR VPWR U$$1034/A sky130_fd_sc_hd__a22o_1
XU$$1044 U$$1044/A U$$1090/B VGND VGND VPWR VPWR U$$1044/X sky130_fd_sc_hd__xor2_1
XFILLER_56_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1055 U$$3245/B1 U$$997/A2 U$$3112/A1 U$$997/B2 VGND VGND VPWR VPWR U$$1056/A sky130_fd_sc_hd__a22o_1
XFILLER_188_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1066 U$$1066/A U$$1078/B VGND VGND VPWR VPWR U$$1066/X sky130_fd_sc_hd__xor2_1
XFILLER_31_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1077 U$$940/A1 U$$1093/A2 U$$940/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1078/A sky130_fd_sc_hd__a22o_1
XU$$1088 U$$1088/A U$$1090/B VGND VGND VPWR VPWR U$$1088/X sky130_fd_sc_hd__xor2_1
XU$$1099 _633_/Q U$$1099/B VGND VGND VPWR VPWR U$$1099/X sky130_fd_sc_hd__and2_1
XFILLER_143_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_110_0 dadda_fa_7_110_0/A dadda_fa_7_110_0/B dadda_fa_7_110_0/CIN VGND
+ VGND VPWR VPWR _535_/D _406_/D sky130_fd_sc_hd__fa_1
XFILLER_192_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_640 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_98_2 U$$3129/X U$$3262/X U$$3395/X VGND VGND VPWR VPWR dadda_fa_3_99_1/B
+ dadda_fa_3_98_3/A sky130_fd_sc_hd__fa_1
XFILLER_176_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_75_1 dadda_fa_5_75_1/A dadda_fa_5_75_1/B dadda_fa_5_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_76_0/B dadda_fa_7_75_0/A sky130_fd_sc_hd__fa_1
XFILLER_137_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1069 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_68_0 dadda_fa_5_68_0/A dadda_fa_5_68_0/B dadda_fa_5_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_69_0/A dadda_fa_6_68_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_8 dadda_fa_1_67_8/A dadda_fa_1_67_8/B dadda_fa_1_67_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_3/A dadda_fa_3_67_0/A sky130_fd_sc_hd__fa_2
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_7_0 dadda_fa_6_7_0/A dadda_fa_6_7_0/B dadda_fa_6_7_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_8_0/B dadda_fa_7_7_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_35_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2290 U$$3521/B1 U$$2326/A2 U$$3386/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2291/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_93_1 U$$2454/X U$$2587/X U$$2720/X VGND VGND VPWR VPWR dadda_fa_2_94_5/B
+ dadda_fa_3_93_0/A sky130_fd_sc_hd__fa_1
XFILLER_162_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_70_0 dadda_fa_4_70_0/A dadda_fa_4_70_0/B dadda_fa_4_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/A dadda_fa_5_70_1/A sky130_fd_sc_hd__fa_1
XFILLER_162_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_86_0 dadda_fa_1_86_0/A U$$1642/X U$$1775/X VGND VGND VPWR VPWR dadda_fa_2_87_2/CIN
+ dadda_fa_2_86_4/B sky130_fd_sc_hd__fa_2
XFILLER_49_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_2_106_1 U$$3278/X U$$3411/X VGND VGND VPWR VPWR dadda_fa_3_107_3/CIN dadda_fa_4_106_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$230 final_adder.U$$725/A final_adder.U$$724/A VGND VGND VPWR VPWR
+ final_adder.U$$306/A sky130_fd_sc_hd__and2_1
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3908 U$$4045/A1 U$$3840/X U$$4456/B1 U$$3841/X VGND VGND VPWR VPWR U$$3909/A sky130_fd_sc_hd__a22o_1
X_601_ _613_/CLK _601_/D VGND VGND VPWR VPWR _601_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3919 U$$3919/A U$$3935/B VGND VGND VPWR VPWR U$$3919/X sky130_fd_sc_hd__xor2_1
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$241 final_adder.U$$735/A final_adder.U$$607/B1 final_adder.U$$241/B1
+ VGND VGND VPWR VPWR final_adder.U$$241/X sky130_fd_sc_hd__a21o_1
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$252 final_adder.U$$747/A final_adder.U$$746/A VGND VGND VPWR VPWR
+ final_adder.U$$252/X sky130_fd_sc_hd__and2_1
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$263 final_adder.U$$262/A final_adder.U$$141/X final_adder.U$$143/X
+ VGND VGND VPWR VPWR final_adder.U$$263/X sky130_fd_sc_hd__a21o_1
XU$$102 U$$648/B1 U$$118/A2 U$$650/B1 U$$118/B2 VGND VGND VPWR VPWR U$$103/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$274 final_adder.U$$274/A final_adder.U$$274/B VGND VGND VPWR VPWR
+ final_adder.U$$328/A sky130_fd_sc_hd__and2_1
XU$$113 U$$113/A U$$117/B VGND VGND VPWR VPWR U$$113/X sky130_fd_sc_hd__xor2_1
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$285 final_adder.U$$284/A final_adder.U$$185/X final_adder.U$$187/X
+ VGND VGND VPWR VPWR final_adder.U$$285/X sky130_fd_sc_hd__a21o_1
XFILLER_205_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$124 U$$946/A1 U$$128/A2 U$$811/A1 U$$128/B2 VGND VGND VPWR VPWR U$$125/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$296 final_adder.U$$296/A final_adder.U$$296/B VGND VGND VPWR VPWR
+ final_adder.U$$340/B sky130_fd_sc_hd__and2_1
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$135 U$$135/A U$$2/A VGND VGND VPWR VPWR U$$135/X sky130_fd_sc_hd__xor2_1
XFILLER_84_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_532_ _534_/CLK _532_/D VGND VGND VPWR VPWR _532_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$146 U$$146/A U$$180/B VGND VGND VPWR VPWR U$$146/X sky130_fd_sc_hd__xor2_1
XFILLER_150_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$157 U$$429/B1 U$$175/A2 U$$707/A1 U$$175/B2 VGND VGND VPWR VPWR U$$158/A sky130_fd_sc_hd__a22o_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$168 U$$168/A U$$196/B VGND VGND VPWR VPWR U$$168/X sky130_fd_sc_hd__xor2_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$179 U$$316/A1 U$$181/A2 U$$44/A1 U$$181/B2 VGND VGND VPWR VPWR U$$180/A sky130_fd_sc_hd__a22o_1
X_463_ _463_/CLK _463_/D VGND VGND VPWR VPWR _463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_394_ _523_/CLK _394_/D VGND VGND VPWR VPWR _394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_448 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_85_0 dadda_fa_6_85_0/A dadda_fa_6_85_0/B dadda_fa_6_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_86_0/B dadda_fa_7_85_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1002 _659_/Q VGND VGND VPWR VPWR U$$3014/A sky130_fd_sc_hd__buf_4
XFILLER_153_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1013 U$$2664/B VGND VGND VPWR VPWR U$$2654/B sky130_fd_sc_hd__buf_6
XFILLER_153_131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1024 _653_/Q VGND VGND VPWR VPWR U$$2531/B sky130_fd_sc_hd__buf_6
Xrepeater1035 U$$2442/B VGND VGND VPWR VPWR U$$2400/B sky130_fd_sc_hd__buf_6
XFILLER_182_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1046 _649_/Q VGND VGND VPWR VPWR U$$2309/B sky130_fd_sc_hd__buf_6
XFILLER_154_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1057 U$$1983/B VGND VGND VPWR VPWR U$$1977/B sky130_fd_sc_hd__buf_6
Xrepeater1068 U$$1884/B VGND VGND VPWR VPWR U$$1852/B sky130_fd_sc_hd__buf_6
XFILLER_5_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1079 U$$1773/B VGND VGND VPWR VPWR U$$1763/B sky130_fd_sc_hd__buf_8
XFILLER_141_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_110 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_861 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$680 U$$817/A1 U$$682/A2 U$$817/B1 U$$682/B2 VGND VGND VPWR VPWR U$$681/A sky130_fd_sc_hd__a22o_1
XU$$691 U$$691/A1 U$$759/A2 U$$828/B1 U$$759/B2 VGND VGND VPWR VPWR U$$692/A sky130_fd_sc_hd__a22o_1
XFILLER_147_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1580 U$$997/A1 VGND VGND VPWR VPWR U$$38/A1 sky130_fd_sc_hd__buf_6
XFILLER_67_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1591 _566_/Q VGND VGND VPWR VPWR U$$3735/A1 sky130_fd_sc_hd__buf_6
XFILLER_99_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_72_6 U$$4407/X input226/X dadda_fa_1_72_6/CIN VGND VGND VPWR VPWR dadda_fa_2_73_2/B
+ dadda_fa_2_72_5/B sky130_fd_sc_hd__fa_1
XFILLER_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_65_5 input218/X dadda_fa_1_65_5/B dadda_fa_1_65_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_66_2/A dadda_fa_2_65_5/A sky130_fd_sc_hd__fa_1
XFILLER_104_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_58_4 U$$3182/X U$$3315/X U$$3448/X VGND VGND VPWR VPWR dadda_fa_2_59_1/CIN
+ dadda_fa_2_58_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_73_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk _634_/CLK VGND VGND VPWR VPWR _637_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_28_2 dadda_fa_4_28_2/A dadda_fa_4_28_2/B dadda_fa_4_28_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/CIN dadda_fa_5_28_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4406 _559_/Q U$$4388/X U$$4408/A1 U$$4430/B2 VGND VGND VPWR VPWR U$$4407/A sky130_fd_sc_hd__a22o_1
XU$$4417 U$$4417/A U$$4417/B VGND VGND VPWR VPWR U$$4417/X sky130_fd_sc_hd__xor2_1
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4428 _570_/Q U$$4388/X U$$4430/A1 U$$4454/B2 VGND VGND VPWR VPWR U$$4429/A sky130_fd_sc_hd__a22o_1
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4439 U$$4439/A U$$4439/B VGND VGND VPWR VPWR U$$4439/X sky130_fd_sc_hd__xor2_1
XU$$3705 U$$3705/A1 U$$3785/A2 U$$3844/A1 U$$3785/B2 VGND VGND VPWR VPWR U$$3706/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3716 U$$3716/A U$$3740/B VGND VGND VPWR VPWR U$$3716/X sky130_fd_sc_hd__xor2_1
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3727 U$$4136/B1 U$$3833/A2 U$$4003/A1 U$$3833/B2 VGND VGND VPWR VPWR U$$3728/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3738 U$$3738/A U$$3740/B VGND VGND VPWR VPWR U$$3738/X sky130_fd_sc_hd__xor2_1
XU$$3749 U$$3884/B1 U$$3785/A2 U$$3751/A1 U$$3785/B2 VGND VGND VPWR VPWR U$$3750/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_2 dadda_fa_3_30_2/A dadda_fa_3_30_2/B dadda_fa_3_30_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_31_1/A dadda_fa_4_30_2/B sky130_fd_sc_hd__fa_2
XFILLER_205_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_320 _237_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_331 _239_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_342 U$$229/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_3_23_1 U$$718/X U$$851/X U$$984/X VGND VGND VPWR VPWR dadda_fa_4_24_0/CIN
+ dadda_fa_4_23_2/A sky130_fd_sc_hd__fa_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_515_ _515_/CLK _515_/D VGND VGND VPWR VPWR _515_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_353 U$$4440/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_364 _623_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_16_0 U$$39/X U$$172/X U$$305/X VGND VGND VPWR VPWR dadda_fa_4_17_1/CIN
+ dadda_fa_4_16_2/B sky130_fd_sc_hd__fa_1
XFILLER_61_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_375 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_386 _622_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_446_ _448_/CLK _446_/D VGND VGND VPWR VPWR _446_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_377_ _507_/CLK _377_/D VGND VGND VPWR VPWR _377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1041 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_82_5 dadda_fa_2_82_5/A dadda_fa_2_82_5/B dadda_fa_2_82_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_2/A dadda_fa_4_82_0/A sky130_fd_sc_hd__fa_2
XFILLER_126_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1039 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_75_4 dadda_fa_2_75_4/A dadda_fa_2_75_4/B dadda_fa_2_75_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/CIN dadda_fa_3_75_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_68_3 dadda_fa_2_68_3/A dadda_fa_2_68_3/B dadda_fa_2_68_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/B dadda_fa_3_68_3/B sky130_fd_sc_hd__fa_1
XFILLER_56_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_38_1 dadda_fa_5_38_1/A dadda_fa_5_38_1/B dadda_fa_5_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_39_0/B dadda_fa_7_38_0/A sky130_fd_sc_hd__fa_2
XFILLER_37_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_75_clk _628_/CLK VGND VGND VPWR VPWR _534_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_1086 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_112_1 dadda_fa_5_112_1/A dadda_fa_5_112_1/B dadda_fa_5_112_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_113_0/B dadda_fa_7_112_0/A sky130_fd_sc_hd__fa_1
XFILLER_192_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_105_0 dadda_fa_5_105_0/A dadda_fa_5_105_0/B dadda_fa_5_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_106_0/A dadda_fa_6_105_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_665 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_315 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_70_3 U$$3472/X U$$3605/X U$$3738/X VGND VGND VPWR VPWR dadda_fa_2_71_1/B
+ dadda_fa_2_70_4/B sky130_fd_sc_hd__fa_1
XFILLER_86_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1092 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_2 U$$3192/X U$$3325/X U$$3458/X VGND VGND VPWR VPWR dadda_fa_2_64_1/A
+ dadda_fa_2_63_4/A sky130_fd_sc_hd__fa_1
XFILLER_115_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_40_1 dadda_fa_4_40_1/A dadda_fa_4_40_1/B dadda_fa_4_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/B dadda_fa_5_40_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_56_1 U$$1582/X U$$1715/X U$$1848/X VGND VGND VPWR VPWR dadda_fa_2_57_0/CIN
+ dadda_fa_2_56_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_33_0 dadda_fa_4_33_0/A dadda_fa_4_33_0/B dadda_fa_4_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/A dadda_fa_5_33_1/A sky130_fd_sc_hd__fa_1
XFILLER_83_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_49_0 U$$105/X U$$238/X U$$371/X VGND VGND VPWR VPWR dadda_fa_2_50_0/CIN
+ dadda_fa_2_49_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_300_ _431_/CLK _300_/D VGND VGND VPWR VPWR _300_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_231_ _353_/CLK _231_/D VGND VGND VPWR VPWR _231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_390 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_85_3 dadda_fa_3_85_3/A dadda_fa_3_85_3/B dadda_fa_3_85_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_1/B dadda_fa_4_85_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_191_590 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_78_2 dadda_fa_3_78_2/A dadda_fa_3_78_2/B dadda_fa_3_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_1/A dadda_fa_4_78_2/B sky130_fd_sc_hd__fa_1
XFILLER_152_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_48_0 dadda_fa_6_48_0/A dadda_fa_6_48_0/B dadda_fa_6_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_49_0/B dadda_fa_7_48_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_211_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4203 U$$4203/A U$$4203/B VGND VGND VPWR VPWR U$$4203/X sky130_fd_sc_hd__xor2_1
XU$$4214 U$$4214/A1 U$$4226/A2 U$$4353/A1 U$$4226/B2 VGND VGND VPWR VPWR U$$4215/A
+ sky130_fd_sc_hd__a22o_1
XU$$4225 U$$4225/A U$$4239/B VGND VGND VPWR VPWR U$$4225/X sky130_fd_sc_hd__xor2_1
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4236 U$$4236/A1 U$$4238/A2 U$$4238/A1 U$$4238/B2 VGND VGND VPWR VPWR U$$4237/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3502 U$$3502/A U$$3506/B VGND VGND VPWR VPWR U$$3502/X sky130_fd_sc_hd__xor2_1
XU$$4247 U$$4247/A VGND VGND VPWR VPWR U$$4247/Y sky130_fd_sc_hd__inv_1
XU$$3513 U$$4333/B1 U$$3537/A2 U$$4198/B1 U$$3537/B2 VGND VGND VPWR VPWR U$$3514/A
+ sky130_fd_sc_hd__a22o_1
XU$$4258 U$$4258/A U$$4298/B VGND VGND VPWR VPWR U$$4258/X sky130_fd_sc_hd__xor2_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_clk _535_/CLK VGND VGND VPWR VPWR _598_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$3524 U$$3524/A U$$3538/B VGND VGND VPWR VPWR U$$3524/X sky130_fd_sc_hd__xor2_1
XU$$4269 U$$4269/A1 U$$4297/A2 U$$4408/A1 U$$4297/B2 VGND VGND VPWR VPWR U$$4270/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3535 U$$3807/B1 U$$3537/A2 _604_/Q U$$3537/B2 VGND VGND VPWR VPWR U$$3536/A sky130_fd_sc_hd__a22o_1
XU$$2801 U$$2801/A U$$2839/B VGND VGND VPWR VPWR U$$2801/X sky130_fd_sc_hd__xor2_1
XU$$3546 U$$3546/A U$$3556/B VGND VGND VPWR VPWR U$$3546/X sky130_fd_sc_hd__xor2_1
XU$$3557 U$$4105/A1 U$$3559/A2 U$$4105/B1 U$$3559/B2 VGND VGND VPWR VPWR U$$3558/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2812 U$$4317/B1 U$$2812/A2 U$$3362/A1 U$$2812/B2 VGND VGND VPWR VPWR U$$2813/A
+ sky130_fd_sc_hd__a22o_1
XU$$2823 U$$2823/A U$$2861/B VGND VGND VPWR VPWR U$$2823/X sky130_fd_sc_hd__xor2_1
XU$$3568 U$$3568/A1 U$$3612/A2 U$$3844/A1 U$$3612/B2 VGND VGND VPWR VPWR U$$3569/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_107_2 dadda_fa_4_107_2/A dadda_fa_4_107_2/B dadda_fa_4_107_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/CIN dadda_fa_5_107_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2834 U$$4478/A1 U$$2874/A2 U$$4480/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2835/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3579 U$$3579/A U$$3613/B VGND VGND VPWR VPWR U$$3579/X sky130_fd_sc_hd__xor2_1
XFILLER_179_808 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2845 U$$2845/A U$$2875/B VGND VGND VPWR VPWR U$$2845/X sky130_fd_sc_hd__xor2_1
XU$$2856 U$$2991/B1 U$$2856/A2 U$$2858/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2857/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2867 U$$2867/A _657_/Q VGND VGND VPWR VPWR U$$2867/X sky130_fd_sc_hd__xor2_1
XANTENNA_150 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _183_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2878 _658_/Q VGND VGND VPWR VPWR U$$2880/B sky130_fd_sc_hd__inv_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2889 U$$3024/B1 U$$2929/A2 U$$3163/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2890/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_429_ _431_/CLK _429_/D VGND VGND VPWR VPWR _429_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_80_2 dadda_fa_2_80_2/A dadda_fa_2_80_2/B dadda_fa_2_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/A dadda_fa_3_80_3/A sky130_fd_sc_hd__fa_1
XFILLER_115_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_73_1 dadda_fa_2_73_1/A dadda_fa_2_73_1/B dadda_fa_2_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_0/CIN dadda_fa_3_73_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_50_0 dadda_fa_5_50_0/A dadda_fa_5_50_0/B dadda_fa_5_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_51_0/A dadda_fa_6_50_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_66_0 dadda_fa_2_66_0/A dadda_fa_2_66_0/B dadda_fa_2_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_0/B dadda_fa_3_66_2/B sky130_fd_sc_hd__fa_1
XFILLER_5_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 a[0] VGND VGND VPWR VPWR _616_/D sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_48_clk _369_/CLK VGND VGND VPWR VPWR _379_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_972 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_95_2 dadda_fa_4_95_2/A dadda_fa_4_95_2/B dadda_fa_4_95_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/CIN dadda_fa_5_95_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_88_1 dadda_fa_4_88_1/A dadda_fa_4_88_1/B dadda_fa_4_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/B dadda_fa_5_88_1/B sky130_fd_sc_hd__fa_1
XFILLER_106_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_65_0 dadda_fa_7_65_0/A dadda_fa_7_65_0/B dadda_fa_7_65_0/CIN VGND VGND
+ VPWR VPWR _490_/D _361_/D sky130_fd_sc_hd__fa_1
XFILLER_126_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput360 _246_/Q VGND VGND VPWR VPWR o[78] sky130_fd_sc_hd__buf_2
XFILLER_0_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput371 _256_/Q VGND VGND VPWR VPWR o[88] sky130_fd_sc_hd__buf_2
Xoutput382 _266_/Q VGND VGND VPWR VPWR o[98] sky130_fd_sc_hd__buf_2
XFILLER_86_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$965_1847 VGND VGND VPWR VPWR U$$965_1847/HI U$$965/A1 sky130_fd_sc_hd__conb_1
XFILLER_0_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_clk _479_/CLK VGND VGND VPWR VPWR _485_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2108 U$$2108/A U$$2108/B VGND VGND VPWR VPWR U$$2108/X sky130_fd_sc_hd__xor2_1
XU$$2119 U$$201/A1 U$$2145/A2 U$$3626/B1 U$$2145/B2 VGND VGND VPWR VPWR U$$2120/A
+ sky130_fd_sc_hd__a22o_1
XU$$1407 U$$1407/A U$$1443/B VGND VGND VPWR VPWR U$$1407/X sky130_fd_sc_hd__xor2_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1418 U$$596/A1 U$$1458/A2 U$$596/B1 U$$1458/B2 VGND VGND VPWR VPWR U$$1419/A sky130_fd_sc_hd__a22o_1
XFILLER_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1429 U$$1429/A U$$1429/B VGND VGND VPWR VPWR U$$1429/X sky130_fd_sc_hd__xor2_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_214_ _475_/CLK _214_/D VGND VGND VPWR VPWR _214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1030 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_90_1 dadda_fa_3_90_1/A dadda_fa_3_90_1/B dadda_fa_3_90_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_0/CIN dadda_fa_4_90_2/A sky130_fd_sc_hd__fa_1
XFILLER_87_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_83_0 dadda_fa_3_83_0/A dadda_fa_3_83_0/B dadda_fa_3_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_0/B dadda_fa_4_83_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4000 U$$4000/A U$$4036/B VGND VGND VPWR VPWR U$$4000/X sky130_fd_sc_hd__xor2_1
XU$$4011 U$$4285/A1 U$$4029/A2 U$$4287/A1 U$$4029/B2 VGND VGND VPWR VPWR U$$4012/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4022 U$$4022/A U$$4044/B VGND VGND VPWR VPWR U$$4022/X sky130_fd_sc_hd__xor2_1
XU$$4033 U$$4168/B1 U$$4035/A2 U$$4035/A1 U$$4081/B2 VGND VGND VPWR VPWR U$$4034/A
+ sky130_fd_sc_hd__a22o_1
XU$$4044 U$$4044/A U$$4044/B VGND VGND VPWR VPWR U$$4044/X sky130_fd_sc_hd__xor2_1
XU$$4055 U$$4466/A1 U$$4061/A2 _590_/Q U$$4061/B2 VGND VGND VPWR VPWR U$$4056/A sky130_fd_sc_hd__a22o_1
XU$$3310 U$$3310/A1 U$$3320/A2 U$$981/B1 U$$3320/B2 VGND VGND VPWR VPWR U$$3311/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4066 U$$4066/A U$$4070/B VGND VGND VPWR VPWR U$$4066/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_0 U$$4354/X U$$4487/X input143/X VGND VGND VPWR VPWR dadda_fa_5_113_0/A
+ dadda_fa_5_112_1/A sky130_fd_sc_hd__fa_1
XFILLER_47_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3321 U$$3321/A U$$3343/B VGND VGND VPWR VPWR U$$3321/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_45_5 dadda_fa_2_45_5/A dadda_fa_2_45_5/B dadda_fa_2_45_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_2/A dadda_fa_4_45_0/A sky130_fd_sc_hd__fa_2
XU$$3332 _570_/Q U$$3368/A2 U$$4430/A1 U$$3368/B2 VGND VGND VPWR VPWR U$$3333/A sky130_fd_sc_hd__a22o_1
XU$$4077 U$$4351/A1 U$$4095/A2 U$$4353/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4078/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3343 U$$3343/A U$$3343/B VGND VGND VPWR VPWR U$$3343/X sky130_fd_sc_hd__xor2_1
XU$$4088 U$$4088/A U$$4109/A VGND VGND VPWR VPWR U$$4088/X sky130_fd_sc_hd__xor2_1
XU$$3354 U$$4450/A1 U$$3404/A2 U$$3354/B1 U$$3404/B2 VGND VGND VPWR VPWR U$$3355/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_38_4 U$$2698/B input188/X dadda_fa_2_38_4/CIN VGND VGND VPWR VPWR dadda_fa_3_39_1/CIN
+ dadda_fa_3_38_3/CIN sky130_fd_sc_hd__fa_1
XU$$4099 U$$4236/A1 U$$4107/A2 U$$4238/A1 U$$4105/B2 VGND VGND VPWR VPWR U$$4100/A
+ sky130_fd_sc_hd__a22o_1
XU$$2620 U$$2620/A U$$2664/B VGND VGND VPWR VPWR U$$2620/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3365 U$$3365/A U$$3407/B VGND VGND VPWR VPWR U$$3365/X sky130_fd_sc_hd__xor2_1
XU$$2631 U$$4273/B1 U$$2697/A2 U$$4140/A1 U$$2697/B2 VGND VGND VPWR VPWR U$$2632/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3376 U$$4472/A1 U$$3408/A2 U$$4472/B1 U$$3408/B2 VGND VGND VPWR VPWR U$$3377/A
+ sky130_fd_sc_hd__a22o_1
XU$$2642 U$$2642/A U$$2688/B VGND VGND VPWR VPWR U$$2642/X sky130_fd_sc_hd__xor2_1
XU$$3387 U$$3387/A U$$3397/B VGND VGND VPWR VPWR U$$3387/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2653 U$$733/B1 U$$2653/A2 U$$3475/B1 U$$2653/B2 VGND VGND VPWR VPWR U$$2654/A
+ sky130_fd_sc_hd__a22o_1
XU$$3398 _603_/Q U$$3402/A2 _604_/Q U$$3402/B2 VGND VGND VPWR VPWR U$$3399/A sky130_fd_sc_hd__a22o_1
XFILLER_146_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2664 U$$2664/A U$$2664/B VGND VGND VPWR VPWR U$$2664/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1930 U$$2613/B1 U$$1956/A2 U$$2754/A1 U$$1956/B2 VGND VGND VPWR VPWR U$$1931/A
+ sky130_fd_sc_hd__a22o_1
XU$$2675 U$$4045/A1 U$$2707/A2 U$$3362/A1 U$$2707/B2 VGND VGND VPWR VPWR U$$2676/A
+ sky130_fd_sc_hd__a22o_1
XU$$2686 U$$2686/A U$$2688/B VGND VGND VPWR VPWR U$$2686/X sky130_fd_sc_hd__xor2_1
XU$$1941 U$$1941/A U$$1977/B VGND VGND VPWR VPWR U$$1941/X sky130_fd_sc_hd__xor2_1
XU$$1952 U$$3320/B1 U$$1956/A2 U$$3735/A1 U$$1956/B2 VGND VGND VPWR VPWR U$$1953/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2697 U$$368/A1 U$$2697/A2 U$$3932/A1 U$$2697/B2 VGND VGND VPWR VPWR U$$2698/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1963 U$$1963/A U$$2011/B VGND VGND VPWR VPWR U$$1963/X sky130_fd_sc_hd__xor2_1
XU$$1974 U$$3618/A1 U$$1976/A2 U$$1976/A1 U$$1976/B2 VGND VGND VPWR VPWR U$$1975/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1985 U$$1985/A U$$2011/B VGND VGND VPWR VPWR U$$1985/X sky130_fd_sc_hd__xor2_1
XU$$1996 U$$624/B1 U$$1922/X U$$491/A1 U$$1923/X VGND VGND VPWR VPWR U$$1997/A sky130_fd_sc_hd__a22o_1
XFILLER_30_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_98_0 dadda_fa_5_98_0/A dadda_fa_5_98_0/B dadda_fa_5_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_99_0/A dadda_fa_6_98_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_590 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$615 final_adder.U$$742/A final_adder.U$$742/B final_adder.U$$615/B1
+ VGND VGND VPWR VPWR final_adder.U$$743/B sky130_fd_sc_hd__a21o_1
XFILLER_69_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$626 final_adder.U$$626/A final_adder.U$$626/B VGND VGND VPWR VPWR
+ _172_/D sky130_fd_sc_hd__xor2_1
Xrepeater830 U$$1923/X VGND VGND VPWR VPWR U$$2040/B2 sky130_fd_sc_hd__buf_8
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater841 U$$1718/B2 VGND VGND VPWR VPWR U$$1710/B2 sky130_fd_sc_hd__buf_6
XFILLER_56_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$637 final_adder.U$$637/A final_adder.U$$637/B VGND VGND VPWR VPWR
+ _183_/D sky130_fd_sc_hd__xor2_4
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater852 U$$1635/B2 VGND VGND VPWR VPWR U$$1627/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$648 final_adder.U$$648/A final_adder.U$$648/B VGND VGND VPWR VPWR
+ _194_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$659 final_adder.U$$659/A final_adder.U$$659/B VGND VGND VPWR VPWR
+ _205_/D sky130_fd_sc_hd__xor2_1
XFILLER_45_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater863 U$$142/X VGND VGND VPWR VPWR U$$263/B2 sky130_fd_sc_hd__buf_4
XFILLER_84_555 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$509 U$$781/B1 U$$517/A2 U$$648/A1 U$$517/B2 VGND VGND VPWR VPWR U$$510/A sky130_fd_sc_hd__a22o_1
Xrepeater874 U$$1291/B2 VGND VGND VPWR VPWR U$$1295/B2 sky130_fd_sc_hd__buf_4
XFILLER_38_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater885 U$$1230/B2 VGND VGND VPWR VPWR U$$1224/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_56_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater896 U$$4438/B2 VGND VGND VPWR VPWR U$$4430/B2 sky130_fd_sc_hd__buf_4
XFILLER_112_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$70 U$$70/A1 U$$84/A2 U$$72/A1 U$$84/B2 VGND VGND VPWR VPWR U$$71/A sky130_fd_sc_hd__a22o_1
XU$$81 U$$81/A U$$81/B VGND VGND VPWR VPWR U$$81/X sky130_fd_sc_hd__xor2_1
XFILLER_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$92 U$$92/A1 U$$98/A2 U$$94/A1 U$$98/B2 VGND VGND VPWR VPWR U$$93/A sky130_fd_sc_hd__a22o_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_496 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_50 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_61 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_94 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1409 U$$4466/A1 VGND VGND VPWR VPWR U$$3779/B1 sky130_fd_sc_hd__buf_4
XFILLER_193_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_730 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_107_1 U$$3812/X U$$3945/X U$$4078/X VGND VGND VPWR VPWR dadda_fa_4_108_0/CIN
+ dadda_fa_4_107_2/A sky130_fd_sc_hd__fa_1
XFILLER_108_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1004 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_48_3 dadda_fa_3_48_3/A dadda_fa_3_48_3/B dadda_fa_3_48_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_1/B dadda_fa_4_48_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1059 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1204 U$$930/A1 U$$1100/X U$$932/A1 U$$1101/X VGND VGND VPWR VPWR U$$1205/A sky130_fd_sc_hd__a22o_1
XFILLER_90_558 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1215 U$$1215/A U$$1225/B VGND VGND VPWR VPWR U$$1215/X sky130_fd_sc_hd__xor2_1
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1226 U$$2459/A1 U$$1230/A2 U$$954/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1227/A
+ sky130_fd_sc_hd__a22o_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1237 U$$1235/Y _634_/Q _633_/Q U$$1236/X U$$1233/Y VGND VGND VPWR VPWR U$$1237/X
+ sky130_fd_sc_hd__a32o_4
XU$$1248 U$$1248/A U$$1296/B VGND VGND VPWR VPWR U$$1248/X sky130_fd_sc_hd__xor2_1
XFILLER_204_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1259 U$$435/B1 U$$1323/A2 U$$302/A1 U$$1323/B2 VGND VGND VPWR VPWR U$$1260/A sky130_fd_sc_hd__a22o_1
XFILLER_141_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_50_3 dadda_fa_2_50_3/A dadda_fa_2_50_3/B dadda_fa_2_50_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/B dadda_fa_3_50_3/B sky130_fd_sc_hd__fa_1
XFILLER_38_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4485_1821 VGND VGND VPWR VPWR U$$4485_1821/HI U$$4485/B sky130_fd_sc_hd__conb_1
XFILLER_39_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_43_2 U$$2753/X U$$2886/X input194/X VGND VGND VPWR VPWR dadda_fa_3_44_1/A
+ dadda_fa_3_43_3/A sky130_fd_sc_hd__fa_1
XFILLER_26_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3140 U$$3412/B1 U$$3144/A2 U$$3551/B1 U$$3144/B2 VGND VGND VPWR VPWR U$$3141/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3151 _661_/Q VGND VGND VPWR VPWR U$$3151/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_5_20_1 dadda_fa_5_20_1/A dadda_fa_5_20_1/B dadda_fa_5_20_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_21_0/B dadda_fa_7_20_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_36_1 U$$1143/X U$$1276/X U$$1409/X VGND VGND VPWR VPWR dadda_fa_3_37_0/CIN
+ dadda_fa_3_36_2/CIN sky130_fd_sc_hd__fa_1
XU$$3162 U$$3162/A U$$3208/B VGND VGND VPWR VPWR U$$3162/X sky130_fd_sc_hd__xor2_1
XFILLER_207_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3173 U$$3310/A1 U$$3215/A2 U$$3175/A1 U$$3215/B2 VGND VGND VPWR VPWR U$$3174/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_13_0 dadda_fa_5_13_0/A dadda_fa_5_13_0/B dadda_fa_5_13_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_14_0/A dadda_fa_6_13_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_81_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3184 U$$3184/A U$$3208/B VGND VGND VPWR VPWR U$$3184/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2450 U$$2450/A U$$2465/A VGND VGND VPWR VPWR U$$2450/X sky130_fd_sc_hd__xor2_1
XU$$3195 U$$4291/A1 U$$3235/A2 U$$4430/A1 U$$3235/B2 VGND VGND VPWR VPWR U$$3196/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2461 _614_/Q U$$2463/A2 _615_/Q U$$2463/B2 VGND VGND VPWR VPWR U$$2462/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_29_0 U$$65/X U$$198/X U$$331/X VGND VGND VPWR VPWR dadda_fa_3_30_1/B dadda_fa_3_29_3/A
+ sky130_fd_sc_hd__fa_1
XFILLER_34_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2472 U$$2472/A1 U$$2550/A2 U$$2611/A1 U$$2550/B2 VGND VGND VPWR VPWR U$$2473/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2483 U$$2483/A U$$2531/B VGND VGND VPWR VPWR U$$2483/X sky130_fd_sc_hd__xor2_1
XU$$2494 U$$987/A1 U$$2516/A2 U$$2494/B1 U$$2516/B2 VGND VGND VPWR VPWR U$$2495/A
+ sky130_fd_sc_hd__a22o_1
XU$$1760 U$$251/B1 U$$1762/A2 U$$253/B1 U$$1762/B2 VGND VGND VPWR VPWR U$$1761/A sky130_fd_sc_hd__a22o_1
XFILLER_179_468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1771 U$$1771/A U$$1773/B VGND VGND VPWR VPWR U$$1771/X sky130_fd_sc_hd__xor2_1
XU$$1782 _642_/Q VGND VGND VPWR VPWR U$$1784/B sky130_fd_sc_hd__inv_1
XU$$1793 U$$971/A1 U$$1859/A2 U$$2754/A1 U$$1859/B2 VGND VGND VPWR VPWR U$$1794/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_803 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput70 b[14] VGND VGND VPWR VPWR _566_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput81 b[24] VGND VGND VPWR VPWR _576_/D sky130_fd_sc_hd__clkbuf_1
Xinput92 b[34] VGND VGND VPWR VPWR _586_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_58_2 dadda_fa_4_58_2/A dadda_fa_4_58_2/B dadda_fa_4_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/CIN dadda_fa_5_58_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$401 final_adder.U$$364/B final_adder.U$$718/B final_adder.U$$345/X
+ VGND VGND VPWR VPWR final_adder.U$$726/B sky130_fd_sc_hd__a21o_4
XTAP_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$423 final_adder.U$$340/B final_adder.U$$702/B final_adder.U$$297/X
+ VGND VGND VPWR VPWR final_adder.U$$706/B sky130_fd_sc_hd__a21o_1
XTAP_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$445 final_adder.U$$268/B final_adder.U$$646/B final_adder.U$$153/X
+ VGND VGND VPWR VPWR final_adder.U$$648/B sky130_fd_sc_hd__a21o_1
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater660 U$$795/B2 VGND VGND VPWR VPWR U$$725/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_7_28_0 dadda_fa_7_28_0/A dadda_fa_7_28_0/B dadda_fa_7_28_0/CIN VGND VGND
+ VPWR VPWR _453_/D _324_/D sky130_fd_sc_hd__fa_1
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater671 U$$553/X VGND VGND VPWR VPWR U$$670/B2 sky130_fd_sc_hd__buf_4
XU$$306 U$$991/A1 U$$308/A2 U$$34/A1 U$$308/B2 VGND VGND VPWR VPWR U$$307/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$467 final_adder.U$$290/B final_adder.U$$690/B final_adder.U$$197/X
+ VGND VGND VPWR VPWR final_adder.U$$692/B sky130_fd_sc_hd__a21o_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$317 U$$317/A U$$351/B VGND VGND VPWR VPWR U$$317/X sky130_fd_sc_hd__xor2_1
Xrepeater682 U$$499/B2 VGND VGND VPWR VPWR U$$483/B2 sky130_fd_sc_hd__buf_4
Xrepeater693 U$$4202/B2 VGND VGND VPWR VPWR U$$4196/B2 sky130_fd_sc_hd__clkbuf_4
XU$$328 U$$463/B1 U$$334/A2 U$$330/A1 U$$334/B2 VGND VGND VPWR VPWR U$$329/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$489 final_adder.U$$312/B final_adder.U$$734/B final_adder.U$$241/X
+ VGND VGND VPWR VPWR final_adder.U$$736/B sky130_fd_sc_hd__a21o_1
XU$$339 U$$339/A U$$351/B VGND VGND VPWR VPWR U$$339/X sky130_fd_sc_hd__xor2_1
XFILLER_199_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_271 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1206 _614_/Q VGND VGND VPWR VPWR U$$3283/A1 sky130_fd_sc_hd__buf_4
Xrepeater1217 U$$948/B1 VGND VGND VPWR VPWR U$$950/A1 sky130_fd_sc_hd__buf_6
XFILLER_5_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1228 U$$3412/B1 VGND VGND VPWR VPWR U$$4236/A1 sky130_fd_sc_hd__buf_4
XFILLER_107_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1239 _610_/Q VGND VGND VPWR VPWR U$$2999/B1 sky130_fd_sc_hd__buf_6
XFILLER_181_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_60_2 dadda_fa_3_60_2/A dadda_fa_3_60_2/B dadda_fa_3_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_1/A dadda_fa_4_60_2/B sky130_fd_sc_hd__fa_1
XFILLER_110_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_53_1 dadda_fa_3_53_1/A dadda_fa_3_53_1/B dadda_fa_3_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_0/CIN dadda_fa_4_53_2/A sky130_fd_sc_hd__fa_1
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_69_1 U$$810/X U$$943/X U$$1076/X VGND VGND VPWR VPWR dadda_fa_1_70_6/B
+ dadda_fa_1_69_8/A sky130_fd_sc_hd__fa_1
XFILLER_121_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_30_0 dadda_fa_6_30_0/A dadda_fa_6_30_0/B dadda_fa_6_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_31_0/B dadda_fa_7_30_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_46_0 dadda_fa_3_46_0/A dadda_fa_3_46_0/B dadda_fa_3_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_0/B dadda_fa_4_46_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$840 U$$840/A1 U$$860/A2 U$$840/B1 U$$860/B2 VGND VGND VPWR VPWR U$$841/A sky130_fd_sc_hd__a22o_1
X_677_ _679_/CLK _677_/D VGND VGND VPWR VPWR _677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$851 U$$851/A U$$925/B VGND VGND VPWR VPWR U$$851/X sky130_fd_sc_hd__xor2_1
XU$$1001 U$$316/A1 U$$979/A2 U$$44/A1 U$$979/B2 VGND VGND VPWR VPWR U$$1002/A sky130_fd_sc_hd__a22o_1
XU$$862 U$$40/A1 U$$928/A2 U$$42/A1 U$$928/B2 VGND VGND VPWR VPWR U$$863/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1012 U$$1012/A U$$980/B VGND VGND VPWR VPWR U$$1012/X sky130_fd_sc_hd__xor2_1
XFILLER_56_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$873 U$$873/A U$$879/B VGND VGND VPWR VPWR U$$873/X sky130_fd_sc_hd__xor2_1
XU$$884 U$$62/A1 U$$928/A2 U$$64/A1 U$$928/B2 VGND VGND VPWR VPWR U$$885/A sky130_fd_sc_hd__a22o_1
XU$$1023 U$$64/A1 U$$1065/A2 U$$66/A1 U$$1065/B2 VGND VGND VPWR VPWR U$$1024/A sky130_fd_sc_hd__a22o_1
XU$$1034 U$$1034/A U$$1040/B VGND VGND VPWR VPWR U$$1034/X sky130_fd_sc_hd__xor2_1
XFILLER_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$895 U$$895/A U$$897/B VGND VGND VPWR VPWR U$$895/X sky130_fd_sc_hd__xor2_1
XU$$1045 U$$908/A1 U$$1089/A2 U$$910/A1 U$$1089/B2 VGND VGND VPWR VPWR U$$1046/A sky130_fd_sc_hd__a22o_1
XFILLER_56_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1056 U$$1056/A U$$998/B VGND VGND VPWR VPWR U$$1056/X sky130_fd_sc_hd__xor2_1
XFILLER_149_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1067 U$$930/A1 U$$963/X U$$932/A1 U$$964/X VGND VGND VPWR VPWR U$$1068/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1078 U$$1078/A U$$1078/B VGND VGND VPWR VPWR U$$1078/X sky130_fd_sc_hd__xor2_1
XU$$1089 U$$952/A1 U$$1089/A2 U$$954/A1 U$$1089/B2 VGND VGND VPWR VPWR U$$1090/A sky130_fd_sc_hd__a22o_1
XFILLER_176_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_103_0 dadda_fa_7_103_0/A dadda_fa_7_103_0/B dadda_fa_7_103_0/CIN VGND
+ VGND VPWR VPWR _528_/D _399_/D sky130_fd_sc_hd__fa_2
XFILLER_184_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_98_3 U$$3528/X U$$3661/X U$$3794/X VGND VGND VPWR VPWR dadda_fa_3_99_1/CIN
+ dadda_fa_3_98_3/B sky130_fd_sc_hd__fa_1
XFILLER_160_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_68_1 dadda_fa_5_68_1/A dadda_fa_5_68_1/B dadda_fa_5_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_69_0/B dadda_fa_7_68_0/A sky130_fd_sc_hd__fa_1
XFILLER_99_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_107_0 U$$3013/Y U$$3147/X U$$3280/X VGND VGND VPWR VPWR dadda_fa_3_108_3/CIN
+ dadda_fa_4_107_0/A sky130_fd_sc_hd__fa_1
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2280 U$$3650/A1 U$$2298/A2 U$$2830/A1 U$$2298/B2 VGND VGND VPWR VPWR U$$2281/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2291 U$$2291/A U$$2328/A VGND VGND VPWR VPWR U$$2291/X sky130_fd_sc_hd__xor2_1
XFILLER_210_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1590 U$$1590/A U$$1598/B VGND VGND VPWR VPWR U$$1590/X sky130_fd_sc_hd__xor2_1
XFILLER_22_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_70_1 dadda_fa_4_70_1/A dadda_fa_4_70_1/B dadda_fa_4_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/B dadda_fa_5_70_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_86_1 U$$1908/X U$$2041/X U$$2174/X VGND VGND VPWR VPWR dadda_fa_2_87_3/A
+ dadda_fa_2_86_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_63_0 dadda_fa_4_63_0/A dadda_fa_4_63_0/B dadda_fa_4_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/A dadda_fa_5_63_1/A sky130_fd_sc_hd__fa_1
XFILLER_77_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_79_0 U$$1095/Y U$$1229/X U$$1362/X VGND VGND VPWR VPWR dadda_fa_2_80_0/B
+ dadda_fa_2_79_3/B sky130_fd_sc_hd__fa_1
XFILLER_131_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$220 final_adder.U$$715/A final_adder.U$$714/A VGND VGND VPWR VPWR
+ final_adder.U$$302/B sky130_fd_sc_hd__and2_1
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$231 final_adder.U$$725/A final_adder.U$$597/B1 final_adder.U$$231/B1
+ VGND VGND VPWR VPWR final_adder.U$$231/X sky130_fd_sc_hd__a21o_1
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_600_ _613_/CLK _600_/D VGND VGND VPWR VPWR _600_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$242 final_adder.U$$737/A final_adder.U$$736/A VGND VGND VPWR VPWR
+ final_adder.U$$312/A sky130_fd_sc_hd__and2_1
XFILLER_73_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3909 U$$3909/A U$$3943/B VGND VGND VPWR VPWR U$$3909/X sky130_fd_sc_hd__xor2_1
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$253 final_adder.U$$747/A final_adder.U$$619/B1 final_adder.U$$253/B1
+ VGND VGND VPWR VPWR final_adder.U$$253/X sky130_fd_sc_hd__a21o_1
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$264 final_adder.U$$264/A final_adder.U$$264/B VGND VGND VPWR VPWR
+ final_adder.U$$324/B sky130_fd_sc_hd__and2_1
XU$$103 U$$103/A U$$117/B VGND VGND VPWR VPWR U$$103/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$275 final_adder.U$$274/A final_adder.U$$165/X final_adder.U$$167/X
+ VGND VGND VPWR VPWR final_adder.U$$275/X sky130_fd_sc_hd__a21o_1
XFILLER_175_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$114 U$$251/A1 U$$118/A2 U$$251/B1 U$$118/B2 VGND VGND VPWR VPWR U$$115/A sky130_fd_sc_hd__a22o_1
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$286 final_adder.U$$286/A final_adder.U$$286/B VGND VGND VPWR VPWR
+ final_adder.U$$334/A sky130_fd_sc_hd__and2_1
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$125 U$$125/A U$$129/B VGND VGND VPWR VPWR U$$125/X sky130_fd_sc_hd__xor2_1
XFILLER_72_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater490 U$$3408/A2 VGND VGND VPWR VPWR U$$3378/A2 sky130_fd_sc_hd__buf_6
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_531_ _559_/CLK _531_/D VGND VGND VPWR VPWR _531_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$297 final_adder.U$$296/A final_adder.U$$209/X final_adder.U$$211/X
+ VGND VGND VPWR VPWR final_adder.U$$297/X sky130_fd_sc_hd__a21o_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$136 _617_/Q VGND VGND VPWR VPWR U$$136/Y sky130_fd_sc_hd__inv_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$147 U$$8/B1 U$$181/A2 U$$12/A1 U$$181/B2 VGND VGND VPWR VPWR U$$148/A sky130_fd_sc_hd__a22o_1
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$158 U$$158/A U$$190/B VGND VGND VPWR VPWR U$$158/X sky130_fd_sc_hd__xor2_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$169 U$$991/A1 U$$195/A2 U$$34/A1 U$$195/B2 VGND VGND VPWR VPWR U$$170/A sky130_fd_sc_hd__a22o_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_462_ _463_/CLK _462_/D VGND VGND VPWR VPWR _462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_393_ _523_/CLK _393_/D VGND VGND VPWR VPWR _393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1003 _657_/Q VGND VGND VPWR VPWR U$$2827/B sky130_fd_sc_hd__buf_8
XFILLER_127_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1014 U$$2706/B VGND VGND VPWR VPWR U$$2664/B sky130_fd_sc_hd__buf_6
Xrepeater1025 _653_/Q VGND VGND VPWR VPWR U$$2567/B sky130_fd_sc_hd__buf_12
Xdadda_fa_6_78_0 dadda_fa_6_78_0/A dadda_fa_6_78_0/B dadda_fa_6_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_79_0/B dadda_fa_7_78_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_153_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1036 U$$2466/A VGND VGND VPWR VPWR U$$2442/B sky130_fd_sc_hd__buf_6
Xrepeater1047 U$$2136/B VGND VGND VPWR VPWR U$$2130/B sky130_fd_sc_hd__buf_8
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1058 U$$2011/B VGND VGND VPWR VPWR U$$1983/B sky130_fd_sc_hd__buf_6
XFILLER_181_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1069 U$$1874/B VGND VGND VPWR VPWR U$$1884/B sky130_fd_sc_hd__buf_8
XFILLER_141_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_124_0_1872 VGND VGND VPWR VPWR dadda_fa_5_124_0/A dadda_fa_5_124_0_1872/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_49_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$670 U$$805/B1 U$$552/X U$$944/B1 U$$670/B2 VGND VGND VPWR VPWR U$$671/A sky130_fd_sc_hd__a22o_1
XFILLER_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$681 U$$681/A U$$684/A VGND VGND VPWR VPWR U$$681/X sky130_fd_sc_hd__xor2_1
XFILLER_211_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_399 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$692 U$$692/A U$$760/B VGND VGND VPWR VPWR U$$692/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_80_0 dadda_fa_5_80_0/A dadda_fa_5_80_0/B dadda_fa_5_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_81_0/A dadda_fa_6_80_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_96_0 U$$2460/X U$$2593/X U$$2726/X VGND VGND VPWR VPWR dadda_fa_3_97_0/B
+ dadda_fa_3_96_2/B sky130_fd_sc_hd__fa_1
XFILLER_172_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1570 _569_/Q VGND VGND VPWR VPWR U$$2508/A1 sky130_fd_sc_hd__buf_4
XFILLER_160_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1581 U$$3187/B1 VGND VGND VPWR VPWR U$$997/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_193_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1592 _566_/Q VGND VGND VPWR VPWR U$$310/A1 sky130_fd_sc_hd__buf_8
XFILLER_98_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_72_7 dadda_fa_1_72_7/A dadda_fa_1_72_7/B dadda_fa_1_72_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_73_2/CIN dadda_fa_2_72_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_65_6 dadda_fa_1_65_6/A dadda_fa_1_65_6/B dadda_fa_1_65_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_2/B dadda_fa_2_65_5/B sky130_fd_sc_hd__fa_1
XFILLER_100_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_58_5 U$$3581/X U$$3714/X U$$3847/X VGND VGND VPWR VPWR dadda_fa_2_59_2/A
+ dadda_fa_2_58_5/A sky130_fd_sc_hd__fa_1
XFILLER_104_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_95_0 dadda_fa_7_95_0/A dadda_fa_7_95_0/B dadda_fa_7_95_0/CIN VGND VGND
+ VPWR VPWR _520_/D _391_/D sky130_fd_sc_hd__fa_1
XFILLER_22_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_750 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4407 U$$4407/A U$$4407/B VGND VGND VPWR VPWR U$$4407/X sky130_fd_sc_hd__xor2_1
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4418 U$$4418/A1 U$$4388/X U$$4418/B1 U$$4430/B2 VGND VGND VPWR VPWR U$$4419/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4429 U$$4429/A U$$4429/B VGND VGND VPWR VPWR U$$4429/X sky130_fd_sc_hd__xor2_1
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_110_0 dadda_fa_6_110_0/A dadda_fa_6_110_0/B dadda_fa_6_110_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_111_0/B dadda_fa_7_110_0/CIN sky130_fd_sc_hd__fa_1
XU$$3706 U$$3706/A U$$3760/B VGND VGND VPWR VPWR U$$3706/X sky130_fd_sc_hd__xor2_1
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3717 _557_/Q U$$3769/A2 U$$3717/B1 U$$3769/B2 VGND VGND VPWR VPWR U$$3718/A sky130_fd_sc_hd__a22o_1
XFILLER_92_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3728 U$$3728/A U$$3832/B VGND VGND VPWR VPWR U$$3728/X sky130_fd_sc_hd__xor2_1
XU$$3739 U$$451/A1 U$$3743/A2 U$$3876/B1 U$$3743/B2 VGND VGND VPWR VPWR U$$3740/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_3 dadda_fa_3_30_3/A dadda_fa_3_30_3/B dadda_fa_3_30_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_31_1/B dadda_fa_4_30_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_310 _236_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 _238_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_23_2 U$$1117/X U$$1250/X U$$1383/X VGND VGND VPWR VPWR dadda_fa_4_24_1/A
+ dadda_fa_4_23_2/B sky130_fd_sc_hd__fa_1
XANTENNA_332 _239_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_514_ _514_/CLK _514_/D VGND VGND VPWR VPWR _514_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_343 U$$229/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_354 U$$3753/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_365 U$$2040/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_376 _634_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_387 U$$1428/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_445_ _445_/CLK _445_/D VGND VGND VPWR VPWR _445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ _507_/CLK _376_/D VGND VGND VPWR VPWR _376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_75_5 dadda_fa_2_75_5/A dadda_fa_2_75_5/B dadda_fa_2_75_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_2/A dadda_fa_4_75_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_4_118_0_1870 VGND VGND VPWR VPWR dadda_fa_4_118_0/A dadda_fa_4_118_0_1870/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_69_915 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_68_4 dadda_fa_2_68_4/A dadda_fa_2_68_4/B dadda_fa_2_68_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/CIN dadda_fa_3_68_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_420 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_599 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_105_1 dadda_fa_5_105_1/A dadda_fa_5_105_1/B dadda_fa_5_105_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_106_0/B dadda_fa_7_105_0/A sky130_fd_sc_hd__fa_1
XFILLER_173_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_414 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_70_4 U$$3871/X U$$4004/X U$$4137/X VGND VGND VPWR VPWR dadda_fa_2_71_1/CIN
+ dadda_fa_2_70_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_119_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_3 U$$3591/X U$$3724/X U$$3857/X VGND VGND VPWR VPWR dadda_fa_2_64_1/B
+ dadda_fa_2_63_4/B sky130_fd_sc_hd__fa_1
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_40_2 dadda_fa_4_40_2/A dadda_fa_4_40_2/B dadda_fa_4_40_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/CIN dadda_fa_5_40_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_56_2 U$$1981/X U$$2114/X U$$2247/X VGND VGND VPWR VPWR dadda_fa_2_57_1/A
+ dadda_fa_2_56_4/A sky130_fd_sc_hd__fa_1
XFILLER_27_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_33_1 dadda_fa_4_33_1/A dadda_fa_4_33_1/B dadda_fa_4_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/B dadda_fa_5_33_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_49_1 U$$504/X U$$637/X U$$770/X VGND VGND VPWR VPWR dadda_fa_2_50_1/A
+ dadda_fa_2_49_4/A sky130_fd_sc_hd__fa_1
XFILLER_55_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_10_0 dadda_fa_7_10_0/A dadda_fa_7_10_0/B dadda_fa_7_10_0/CIN VGND VGND
+ VPWR VPWR _435_/D _306_/D sky130_fd_sc_hd__fa_1
XFILLER_54_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_26_0 dadda_fa_4_26_0/A dadda_fa_4_26_0/B dadda_fa_4_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/A dadda_fa_5_26_1/A sky130_fd_sc_hd__fa_1
XFILLER_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_230_ _353_/CLK _230_/D VGND VGND VPWR VPWR _230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_78_3 dadda_fa_3_78_3/A dadda_fa_3_78_3/B dadda_fa_3_78_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_1/B dadda_fa_4_78_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4204 _595_/Q U$$4114/X _596_/Q U$$4115/X VGND VGND VPWR VPWR U$$4205/A sky130_fd_sc_hd__a22o_1
XFILLER_93_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4215 U$$4215/A U$$4215/B VGND VGND VPWR VPWR U$$4215/X sky130_fd_sc_hd__xor2_1
XFILLER_172_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4226 U$$4361/B1 U$$4226/A2 U$$4500/B1 U$$4226/B2 VGND VGND VPWR VPWR U$$4227/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4237 U$$4237/A U$$4239/B VGND VGND VPWR VPWR U$$4237/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_3_15_0 U$$37/X U$$170/X VGND VGND VPWR VPWR dadda_fa_4_16_2/A dadda_ha_3_15_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$3503 U$$3503/A1 U$$3545/A2 U$$3642/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3504/A
+ sky130_fd_sc_hd__a22o_1
XU$$4248 _678_/Q VGND VGND VPWR VPWR U$$4250/B sky130_fd_sc_hd__inv_1
XU$$3514 U$$3514/A U$$3520/B VGND VGND VPWR VPWR U$$3514/X sky130_fd_sc_hd__xor2_1
XU$$4259 U$$4396/A1 U$$4297/A2 U$$4259/B1 U$$4297/B2 VGND VGND VPWR VPWR U$$4260/A
+ sky130_fd_sc_hd__a22o_1
XU$$3525 _598_/Q U$$3531/A2 _599_/Q U$$3531/B2 VGND VGND VPWR VPWR U$$3526/A sky130_fd_sc_hd__a22o_1
XFILLER_92_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3536 U$$3536/A U$$3562/A VGND VGND VPWR VPWR U$$3536/X sky130_fd_sc_hd__xor2_1
XU$$2802 U$$4035/A1 U$$2832/A2 U$$4035/B1 U$$2832/B2 VGND VGND VPWR VPWR U$$2803/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3547 U$$4506/A1 U$$3555/A2 U$$4508/A1 U$$3555/B2 VGND VGND VPWR VPWR U$$3548/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3558 U$$3558/A U$$3561/A VGND VGND VPWR VPWR U$$3558/X sky130_fd_sc_hd__xor2_1
XU$$2813 U$$2813/A U$$2813/B VGND VGND VPWR VPWR U$$2813/X sky130_fd_sc_hd__xor2_1
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2824 U$$3783/A1 U$$2856/A2 U$$4194/B1 U$$2856/B2 VGND VGND VPWR VPWR U$$2825/A
+ sky130_fd_sc_hd__a22o_1
XU$$3569 U$$3569/A U$$3613/B VGND VGND VPWR VPWR U$$3569/X sky130_fd_sc_hd__xor2_1
XFILLER_45_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2835 U$$2835/A U$$2877/A VGND VGND VPWR VPWR U$$2835/X sky130_fd_sc_hd__xor2_1
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2846 U$$3942/A1 U$$2866/A2 U$$2983/B1 U$$2866/B2 VGND VGND VPWR VPWR U$$2847/A
+ sky130_fd_sc_hd__a22o_1
XU$$2857 U$$2857/A U$$2861/B VGND VGND VPWR VPWR U$$2857/X sky130_fd_sc_hd__xor2_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _290_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2868 U$$3551/B1 U$$2874/A2 U$$3281/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2869/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_151 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _183_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2879 U$$3014/A VGND VGND VPWR VPWR U$$2879/Y sky130_fd_sc_hd__inv_1
XANTENNA_173 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_195 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_428_ _428_/CLK _428_/D VGND VGND VPWR VPWR _428_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_359_ _488_/CLK _359_/D VGND VGND VPWR VPWR _359_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_80_3 dadda_fa_2_80_3/A dadda_fa_2_80_3/B dadda_fa_2_80_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/B dadda_fa_3_80_3/B sky130_fd_sc_hd__fa_1
XFILLER_142_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_73_2 dadda_fa_2_73_2/A dadda_fa_2_73_2/B dadda_fa_2_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/A dadda_fa_3_73_3/A sky130_fd_sc_hd__fa_1
XFILLER_155_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_50_1 dadda_fa_5_50_1/A dadda_fa_5_50_1/B dadda_fa_5_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_51_0/B dadda_fa_7_50_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_66_1 dadda_fa_2_66_1/A dadda_fa_2_66_1/B dadda_fa_2_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_0/CIN dadda_fa_3_66_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_1176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4449_1803 VGND VGND VPWR VPWR U$$4449_1803/HI U$$4449/B sky130_fd_sc_hd__conb_1
Xdadda_fa_5_43_0 dadda_fa_5_43_0/A dadda_fa_5_43_0/B dadda_fa_5_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_44_0/A dadda_fa_6_43_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_59_0 dadda_fa_2_59_0/A dadda_fa_2_59_0/B dadda_fa_2_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_0/B dadda_fa_3_59_2/B sky130_fd_sc_hd__fa_1
Xinput2 a[10] VGND VGND VPWR VPWR _626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_859 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$0 _424_/Q _296_/Q VGND VGND VPWR VPWR final_adder.U$$623/B final_adder.U$$622/A
+ sky130_fd_sc_hd__ha_1
XFILLER_192_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_88_2 dadda_fa_4_88_2/A dadda_fa_4_88_2/B dadda_fa_4_88_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/CIN dadda_fa_5_88_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput350 _237_/Q VGND VGND VPWR VPWR o[69] sky130_fd_sc_hd__buf_2
XFILLER_160_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput361 _247_/Q VGND VGND VPWR VPWR o[79] sky130_fd_sc_hd__buf_2
Xdadda_fa_7_58_0 dadda_fa_7_58_0/A dadda_fa_7_58_0/B dadda_fa_7_58_0/CIN VGND VGND
+ VPWR VPWR _483_/D _354_/D sky130_fd_sc_hd__fa_1
XFILLER_133_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput372 _257_/Q VGND VGND VPWR VPWR o[89] sky130_fd_sc_hd__buf_2
XFILLER_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput383 _267_/Q VGND VGND VPWR VPWR o[99] sky130_fd_sc_hd__buf_2
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_0 U$$1991/X U$$2124/X U$$2257/X VGND VGND VPWR VPWR dadda_fa_2_62_0/B
+ dadda_fa_2_61_3/B sky130_fd_sc_hd__fa_1
XFILLER_47_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4389_1772 VGND VGND VPWR VPWR U$$4389_1772/HI U$$4389/B1 sky130_fd_sc_hd__conb_1
XFILLER_90_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2109 U$$3753/A1 U$$2109/A2 U$$3618/A1 U$$2109/B2 VGND VGND VPWR VPWR U$$2110/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1408 U$$2641/A1 U$$1442/A2 U$$2641/B1 U$$1442/B2 VGND VGND VPWR VPWR U$$1409/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1419 U$$1419/A U$$1459/B VGND VGND VPWR VPWR U$$1419/X sky130_fd_sc_hd__xor2_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_213_ _213_/CLK _213_/D VGND VGND VPWR VPWR _213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1001 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_90_2 dadda_fa_3_90_2/A dadda_fa_3_90_2/B dadda_fa_3_90_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_1/A dadda_fa_4_90_2/B sky130_fd_sc_hd__fa_1
XFILLER_137_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_83_1 dadda_fa_3_83_1/A dadda_fa_3_83_1/B dadda_fa_3_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_0/CIN dadda_fa_4_83_2/A sky130_fd_sc_hd__fa_1
XFILLER_83_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_60_0 dadda_fa_6_60_0/A dadda_fa_6_60_0/B dadda_fa_6_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_61_0/B dadda_fa_7_60_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_76_0 dadda_fa_3_76_0/A dadda_fa_3_76_0/B dadda_fa_3_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_0/B dadda_fa_4_76_1/CIN sky130_fd_sc_hd__fa_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4001 U$$4136/B1 U$$4035/A2 U$$4003/A1 U$$4081/B2 VGND VGND VPWR VPWR U$$4002/A
+ sky130_fd_sc_hd__a22o_1
XU$$4012 U$$4012/A U$$4044/B VGND VGND VPWR VPWR U$$4012/X sky130_fd_sc_hd__xor2_1
XU$$4023 U$$4160/A1 U$$4029/A2 _574_/Q U$$4029/B2 VGND VGND VPWR VPWR U$$4024/A sky130_fd_sc_hd__a22o_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4034 U$$4034/A U$$4096/B VGND VGND VPWR VPWR U$$4034/X sky130_fd_sc_hd__xor2_1
XU$$3300 U$$3437/A1 U$$3320/A2 U$$3713/A1 U$$3320/B2 VGND VGND VPWR VPWR U$$3301/A
+ sky130_fd_sc_hd__a22o_1
XU$$4045 U$$4045/A1 U$$4065/A2 U$$4456/B1 U$$4065/B2 VGND VGND VPWR VPWR U$$4046/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3311 U$$3311/A U$$3363/B VGND VGND VPWR VPWR U$$3311/X sky130_fd_sc_hd__xor2_1
XU$$4056 U$$4056/A U$$4058/B VGND VGND VPWR VPWR U$$4056/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_1 dadda_fa_4_112_1/A dadda_fa_4_112_1/B dadda_fa_4_112_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_113_0/B dadda_fa_5_112_1/B sky130_fd_sc_hd__fa_1
XU$$4067 _595_/Q U$$4071/A2 _596_/Q U$$4071/B2 VGND VGND VPWR VPWR U$$4068/A sky130_fd_sc_hd__a22o_1
XFILLER_20_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3322 U$$4007/A1 U$$3368/A2 U$$3735/A1 U$$3368/B2 VGND VGND VPWR VPWR U$$3323/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3333 U$$3333/A U$$3369/B VGND VGND VPWR VPWR U$$3333/X sky130_fd_sc_hd__xor2_1
XU$$4078 U$$4078/A U$$4084/B VGND VGND VPWR VPWR U$$4078/X sky130_fd_sc_hd__xor2_1
XU$$3344 U$$4027/B1 U$$3356/A2 U$$3346/A1 U$$3356/B2 VGND VGND VPWR VPWR U$$3345/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4089 U$$4361/B1 U$$4095/A2 U$$4500/B1 U$$4105/B2 VGND VGND VPWR VPWR U$$4090/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_754 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3355 U$$3355/A U$$3397/B VGND VGND VPWR VPWR U$$3355/X sky130_fd_sc_hd__xor2_1
XU$$2610 U$$2610/A U$$2698/B VGND VGND VPWR VPWR U$$2610/X sky130_fd_sc_hd__xor2_1
XFILLER_93_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2621 U$$2893/B1 U$$2653/A2 U$$3717/B1 U$$2653/B2 VGND VGND VPWR VPWR U$$2622/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_105_0 dadda_fa_4_105_0/A dadda_fa_4_105_0/B dadda_fa_4_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/A dadda_fa_5_105_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_38_5 dadda_fa_2_38_5/A dadda_fa_2_38_5/B dadda_fa_2_38_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_39_2/A dadda_fa_4_38_0/A sky130_fd_sc_hd__fa_2
XFILLER_62_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3366 U$$3503/A1 U$$3418/A2 U$$3642/A1 U$$3418/B2 VGND VGND VPWR VPWR U$$3367/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2632 U$$2632/A U$$2698/B VGND VGND VPWR VPWR U$$2632/X sky130_fd_sc_hd__xor2_1
XU$$3377 U$$3377/A U$$3407/B VGND VGND VPWR VPWR U$$3377/X sky130_fd_sc_hd__xor2_1
XU$$2643 U$$4287/A1 U$$2687/A2 _569_/Q U$$2687/B2 VGND VGND VPWR VPWR U$$2644/A sky130_fd_sc_hd__a22o_1
XU$$3388 _598_/Q U$$3402/A2 U$$3388/B1 U$$3402/B2 VGND VGND VPWR VPWR U$$3389/A sky130_fd_sc_hd__a22o_1
XFILLER_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_943 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3399 U$$3399/A _665_/Q VGND VGND VPWR VPWR U$$3399/X sky130_fd_sc_hd__xor2_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2654 U$$2654/A U$$2654/B VGND VGND VPWR VPWR U$$2654/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2665 U$$4035/A1 U$$2705/A2 U$$4035/B1 U$$2705/B2 VGND VGND VPWR VPWR U$$2666/A
+ sky130_fd_sc_hd__a22o_1
XU$$1920 _645_/Q VGND VGND VPWR VPWR U$$1920/Y sky130_fd_sc_hd__inv_1
XFILLER_55_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1931 U$$1931/A U$$1957/B VGND VGND VPWR VPWR U$$1931/X sky130_fd_sc_hd__xor2_1
XU$$2676 U$$2676/A U$$2708/B VGND VGND VPWR VPWR U$$2676/X sky130_fd_sc_hd__xor2_1
XU$$1942 U$$2077/B1 U$$1982/A2 U$$848/A1 U$$1982/B2 VGND VGND VPWR VPWR U$$1943/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2687 U$$3783/A1 U$$2687/A2 U$$908/A1 U$$2687/B2 VGND VGND VPWR VPWR U$$2688/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1953 U$$1953/A U$$1957/B VGND VGND VPWR VPWR U$$1953/X sky130_fd_sc_hd__xor2_1
XU$$2698 U$$2698/A U$$2698/B VGND VGND VPWR VPWR U$$2698/X sky130_fd_sc_hd__xor2_1
XU$$1964 U$$46/A1 U$$1982/A2 U$$2375/B1 U$$1982/B2 VGND VGND VPWR VPWR U$$1965/A sky130_fd_sc_hd__a22o_1
XU$$1975 U$$1975/A U$$1977/B VGND VGND VPWR VPWR U$$1975/X sky130_fd_sc_hd__xor2_1
XFILLER_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1986 U$$3493/A1 U$$2010/A2 U$$3495/A1 U$$2010/B2 VGND VGND VPWR VPWR U$$1987/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4479_1818 VGND VGND VPWR VPWR U$$4479_1818/HI U$$4479/B sky130_fd_sc_hd__conb_1
XU$$1997 U$$1997/A U$$2003/B VGND VGND VPWR VPWR U$$1997/X sky130_fd_sc_hd__xor2_1
XFILLER_187_694 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_98_1 dadda_fa_5_98_1/A dadda_fa_5_98_1/B dadda_fa_5_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_99_0/B dadda_fa_7_98_0/A sky130_fd_sc_hd__fa_1
XFILLER_174_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$605 final_adder.U$$732/A final_adder.U$$732/B final_adder.U$$605/B1
+ VGND VGND VPWR VPWR final_adder.U$$733/B sky130_fd_sc_hd__a21o_1
Xrepeater820 U$$2060/X VGND VGND VPWR VPWR U$$2169/B2 sky130_fd_sc_hd__buf_4
XFILLER_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$627 final_adder.U$$627/A final_adder.U$$627/B VGND VGND VPWR VPWR
+ _173_/D sky130_fd_sc_hd__xor2_1
XFILLER_29_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_1029 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater831 U$$1786/X VGND VGND VPWR VPWR U$$1859/B2 sky130_fd_sc_hd__buf_6
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$638 final_adder.U$$638/A final_adder.U$$638/B VGND VGND VPWR VPWR
+ _184_/D sky130_fd_sc_hd__xor2_4
Xrepeater842 U$$1768/B2 VGND VGND VPWR VPWR U$$1718/B2 sky130_fd_sc_hd__buf_4
XFILLER_56_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$649 final_adder.U$$649/A final_adder.U$$649/B VGND VGND VPWR VPWR
+ _195_/D sky130_fd_sc_hd__xor2_4
Xrepeater853 U$$1635/B2 VGND VGND VPWR VPWR U$$1587/B2 sky130_fd_sc_hd__buf_6
Xrepeater864 U$$1458/B2 VGND VGND VPWR VPWR U$$1424/B2 sky130_fd_sc_hd__buf_4
Xrepeater875 U$$1323/B2 VGND VGND VPWR VPWR U$$1291/B2 sky130_fd_sc_hd__buf_6
XFILLER_84_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater886 U$$1208/B2 VGND VGND VPWR VPWR U$$1230/B2 sky130_fd_sc_hd__buf_8
Xrepeater897 U$$4389/X VGND VGND VPWR VPWR U$$4438/B2 sky130_fd_sc_hd__buf_6
XFILLER_53_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$60 U$$60/A1 U$$62/A2 U$$62/A1 U$$62/B2 VGND VGND VPWR VPWR U$$61/A sky130_fd_sc_hd__a22o_1
XU$$71 U$$71/A U$$85/B VGND VGND VPWR VPWR U$$71/X sky130_fd_sc_hd__xor2_1
XU$$82 U$$82/A1 U$$84/A2 U$$84/A1 U$$84/B2 VGND VGND VPWR VPWR U$$83/A sky130_fd_sc_hd__a22o_1
XFILLER_198_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$93 U$$93/A U$$93/B VGND VGND VPWR VPWR U$$93/X sky130_fd_sc_hd__xor2_1
XFILLER_72_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4503_1830 VGND VGND VPWR VPWR U$$4503_1830/HI U$$4503/B sky130_fd_sc_hd__conb_1
XFILLER_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_40 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_51 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_62 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_84 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_93_0 dadda_fa_4_93_0/A dadda_fa_4_93_0/B dadda_fa_4_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/A dadda_fa_5_93_1/A sky130_fd_sc_hd__fa_1
XFILLER_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_95 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_336 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_107_2 U$$4211/X U$$4344/X U$$4477/X VGND VGND VPWR VPWR dadda_fa_4_108_1/A
+ dadda_fa_4_107_2/B sky130_fd_sc_hd__fa_1
XFILLER_122_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1205 U$$1205/A _633_/Q VGND VGND VPWR VPWR U$$1205/X sky130_fd_sc_hd__xor2_1
XU$$1216 U$$942/A1 U$$1230/A2 U$$942/B1 U$$1230/B2 VGND VGND VPWR VPWR U$$1217/A sky130_fd_sc_hd__a22o_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1227 U$$1227/A U$$1232/A VGND VGND VPWR VPWR U$$1227/X sky130_fd_sc_hd__xor2_1
XFILLER_16_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1238 U$$1236/B _633_/Q _634_/Q U$$1233/Y VGND VGND VPWR VPWR U$$1238/X sky130_fd_sc_hd__a22o_4
XFILLER_71_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1249 U$$973/B1 U$$1295/A2 U$$429/A1 U$$1295/B2 VGND VGND VPWR VPWR U$$1250/A sky130_fd_sc_hd__a22o_1
XFILLER_102_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_840 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_506 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_50_4 dadda_fa_2_50_4/A dadda_fa_2_50_4/B dadda_fa_2_50_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/CIN dadda_fa_3_50_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_43_3 dadda_fa_2_43_3/A dadda_fa_2_43_3/B dadda_fa_2_43_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_1/B dadda_fa_3_43_3/B sky130_fd_sc_hd__fa_1
XU$$3130 _606_/Q U$$3132/A2 U$$3132/A1 U$$3132/B2 VGND VGND VPWR VPWR U$$3131/A sky130_fd_sc_hd__a22o_1
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3141 U$$3141/A U$$3145/B VGND VGND VPWR VPWR U$$3141/X sky130_fd_sc_hd__xor2_1
XU$$3152 _662_/Q VGND VGND VPWR VPWR U$$3154/B sky130_fd_sc_hd__inv_1
XFILLER_81_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_36_2 U$$1542/X U$$1675/X U$$1808/X VGND VGND VPWR VPWR dadda_fa_3_37_1/A
+ dadda_fa_3_36_3/A sky130_fd_sc_hd__fa_1
XU$$3163 U$$3437/A1 U$$3209/A2 U$$3163/B1 U$$3209/B2 VGND VGND VPWR VPWR U$$3164/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3174 U$$3174/A U$$3218/B VGND VGND VPWR VPWR U$$3174/X sky130_fd_sc_hd__xor2_1
XU$$2440 U$$2440/A U$$2466/A VGND VGND VPWR VPWR U$$2440/X sky130_fd_sc_hd__xor2_1
XU$$3185 U$$3320/B1 U$$3209/A2 U$$856/B1 U$$3209/B2 VGND VGND VPWR VPWR U$$3186/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_13_1 dadda_fa_5_13_1/A dadda_fa_5_13_1/B dadda_ha_4_13_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_14_0/B dadda_fa_7_13_0/A sky130_fd_sc_hd__fa_2
XU$$2451 U$$2586/B1 U$$2451/A2 _610_/Q U$$2451/B2 VGND VGND VPWR VPWR U$$2452/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_29_1 U$$464/X U$$597/X U$$730/X VGND VGND VPWR VPWR dadda_fa_3_30_1/CIN
+ dadda_fa_3_29_3/B sky130_fd_sc_hd__fa_1
XU$$3196 U$$3196/A U$$3236/B VGND VGND VPWR VPWR U$$3196/X sky130_fd_sc_hd__xor2_1
XFILLER_50_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2462 U$$2462/A U$$2462/B VGND VGND VPWR VPWR U$$2462/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2473 U$$2473/A U$$2517/B VGND VGND VPWR VPWR U$$2473/X sky130_fd_sc_hd__xor2_1
XFILLER_34_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2484 U$$2756/B1 U$$2530/A2 U$$840/B1 U$$2530/B2 VGND VGND VPWR VPWR U$$2485/A
+ sky130_fd_sc_hd__a22o_1
XU$$1750 U$$791/A1 U$$1762/A2 U$$517/B1 U$$1762/B2 VGND VGND VPWR VPWR U$$1751/A sky130_fd_sc_hd__a22o_1
XU$$2495 U$$2495/A U$$2541/B VGND VGND VPWR VPWR U$$2495/X sky130_fd_sc_hd__xor2_1
XU$$1761 U$$1761/A U$$1763/B VGND VGND VPWR VPWR U$$1761/X sky130_fd_sc_hd__xor2_1
XFILLER_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1772 U$$950/A1 U$$1778/A2 U$$3418/A1 U$$1778/B2 VGND VGND VPWR VPWR U$$1773/A
+ sky130_fd_sc_hd__a22o_1
XU$$1783 U$$1918/A VGND VGND VPWR VPWR U$$1783/Y sky130_fd_sc_hd__inv_1
XFILLER_188_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1794 U$$1794/A U$$1820/B VGND VGND VPWR VPWR U$$1794/X sky130_fd_sc_hd__xor2_1
XFILLER_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_623 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput60 a[63] VGND VGND VPWR VPWR _679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput71 b[15] VGND VGND VPWR VPWR _567_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput82 b[25] VGND VGND VPWR VPWR _577_/D sky130_fd_sc_hd__clkbuf_1
Xinput93 b[35] VGND VGND VPWR VPWR _587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1010 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1057 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_810 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$413 final_adder.U$$330/B final_adder.U$$662/B final_adder.U$$277/X
+ VGND VGND VPWR VPWR final_adder.U$$666/B sky130_fd_sc_hd__a21o_4
Xfinal_adder.U$$435 final_adder.U$$258/B final_adder.U$$626/B final_adder.U$$133/X
+ VGND VGND VPWR VPWR final_adder.U$$628/B sky130_fd_sc_hd__a21o_1
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater650 U$$896/B2 VGND VGND VPWR VPWR U$$878/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_85_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$457 final_adder.U$$280/B final_adder.U$$670/B final_adder.U$$177/X
+ VGND VGND VPWR VPWR final_adder.U$$672/B sky130_fd_sc_hd__a21o_1
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater661 U$$795/B2 VGND VGND VPWR VPWR U$$759/B2 sky130_fd_sc_hd__buf_6
XFILLER_123_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater672 U$$4333/B2 VGND VGND VPWR VPWR U$$4319/B2 sky130_fd_sc_hd__buf_4
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$307 U$$307/A U$$335/B VGND VGND VPWR VPWR U$$307/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$479 final_adder.U$$302/B final_adder.U$$714/B final_adder.U$$221/X
+ VGND VGND VPWR VPWR final_adder.U$$716/B sky130_fd_sc_hd__a21o_1
Xrepeater683 U$$491/B2 VGND VGND VPWR VPWR U$$499/B2 sky130_fd_sc_hd__buf_6
XFILLER_42_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$318 U$$866/A1 U$$318/A2 U$$866/B1 U$$318/B2 VGND VGND VPWR VPWR U$$319/A sky130_fd_sc_hd__a22o_1
XU$$329 U$$329/A U$$397/B VGND VGND VPWR VPWR U$$329/X sky130_fd_sc_hd__xor2_1
Xrepeater694 U$$4115/X VGND VGND VPWR VPWR U$$4202/B2 sky130_fd_sc_hd__buf_6
XFILLER_84_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1207 _614_/Q VGND VGND VPWR VPWR U$$2459/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_112_0 dadda_fa_3_112_0/A U$$3423/X U$$3556/X VGND VGND VPWR VPWR dadda_fa_4_113_1/B
+ dadda_fa_4_112_2/A sky130_fd_sc_hd__fa_1
XFILLER_10_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1218 _612_/Q VGND VGND VPWR VPWR U$$948/B1 sky130_fd_sc_hd__buf_6
XFILLER_10_1023 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1229 U$$3412/B1 VGND VGND VPWR VPWR U$$4510/A1 sky130_fd_sc_hd__buf_4
XFILLER_107_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_60_3 dadda_fa_3_60_3/A dadda_fa_3_60_3/B dadda_fa_3_60_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_1/B dadda_fa_4_60_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_53_2 dadda_fa_3_53_2/A dadda_fa_3_53_2/B dadda_fa_3_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_1/A dadda_fa_4_53_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_0_69_2 U$$1209/X U$$1342/X U$$1475/X VGND VGND VPWR VPWR dadda_fa_1_70_6/CIN
+ dadda_fa_1_69_8/B sky130_fd_sc_hd__fa_1
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_46_1 dadda_fa_3_46_1/A dadda_fa_3_46_1/B dadda_fa_3_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_0/CIN dadda_fa_4_46_2/A sky130_fd_sc_hd__fa_1
XTAP_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1034 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_23_0 dadda_fa_6_23_0/A dadda_fa_6_23_0/B dadda_fa_6_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_24_0/B dadda_fa_7_23_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_39_0 dadda_fa_3_39_0/A dadda_fa_3_39_0/B dadda_fa_3_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_0/B dadda_fa_4_39_1/CIN sky130_fd_sc_hd__fa_1
XU$$830 U$$967/A1 U$$860/A2 U$$969/A1 U$$860/B2 VGND VGND VPWR VPWR U$$831/A sky130_fd_sc_hd__a22o_1
X_676_ _679_/CLK _676_/D VGND VGND VPWR VPWR _676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$841 U$$841/A U$$859/B VGND VGND VPWR VPWR U$$841/X sky130_fd_sc_hd__xor2_1
XFILLER_169_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$852 U$$30/A1 U$$924/A2 U$$854/A1 U$$924/B2 VGND VGND VPWR VPWR U$$853/A sky130_fd_sc_hd__a22o_1
XU$$1002 U$$1002/A U$$980/B VGND VGND VPWR VPWR U$$1002/X sky130_fd_sc_hd__xor2_1
XFILLER_17_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$863 U$$863/A U$$929/B VGND VGND VPWR VPWR U$$863/X sky130_fd_sc_hd__xor2_1
XU$$874 U$$874/A1 U$$878/A2 U$$876/A1 U$$878/B2 VGND VGND VPWR VPWR U$$875/A sky130_fd_sc_hd__a22o_1
XU$$1013 U$$52/B1 U$$999/A2 U$$467/A1 U$$999/B2 VGND VGND VPWR VPWR U$$1014/A sky130_fd_sc_hd__a22o_1
XU$$1024 U$$1024/A U$$996/B VGND VGND VPWR VPWR U$$1024/X sky130_fd_sc_hd__xor2_1
XU$$885 U$$885/A U$$935/B VGND VGND VPWR VPWR U$$885/X sky130_fd_sc_hd__xor2_1
XFILLER_204_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1035 U$$898/A1 U$$1039/A2 U$$78/A1 U$$1039/B2 VGND VGND VPWR VPWR U$$1036/A sky130_fd_sc_hd__a22o_1
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$896 U$$896/A1 U$$896/A2 U$$896/B1 U$$896/B2 VGND VGND VPWR VPWR U$$897/A sky130_fd_sc_hd__a22o_1
XU$$1046 U$$1046/A U$$1090/B VGND VGND VPWR VPWR U$$1046/X sky130_fd_sc_hd__xor2_1
XFILLER_31_412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1057 U$$98/A1 U$$997/A2 U$$98/B1 U$$997/B2 VGND VGND VPWR VPWR U$$1058/A sky130_fd_sc_hd__a22o_1
XU$$1068 U$$1068/A U$$1078/B VGND VGND VPWR VPWR U$$1068/X sky130_fd_sc_hd__xor2_1
XFILLER_204_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1079 U$$3132/B1 U$$1093/A2 U$$944/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1080/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_98_4 U$$3927/X U$$4060/X U$$4193/X VGND VGND VPWR VPWR dadda_fa_3_99_2/A
+ dadda_fa_3_98_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_41_0 U$$1552/X U$$1685/X U$$1818/X VGND VGND VPWR VPWR dadda_fa_3_42_0/B
+ dadda_fa_3_41_2/B sky130_fd_sc_hd__fa_1
XFILLER_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2270 U$$3503/A1 U$$2274/A2 U$$3642/A1 U$$2274/B2 VGND VGND VPWR VPWR U$$2271/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2281 U$$2281/A U$$2299/B VGND VGND VPWR VPWR U$$2281/X sky130_fd_sc_hd__xor2_1
XU$$2292 U$$3386/B1 U$$2318/A2 U$$785/B1 U$$2318/B2 VGND VGND VPWR VPWR U$$2293/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1580 U$$1580/A U$$1628/B VGND VGND VPWR VPWR U$$1580/X sky130_fd_sc_hd__xor2_1
XFILLER_167_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1591 U$$358/A1 U$$1597/A2 U$$86/A1 U$$1597/B2 VGND VGND VPWR VPWR U$$1592/A sky130_fd_sc_hd__a22o_1
XFILLER_210_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_70_2 dadda_fa_4_70_2/A dadda_fa_4_70_2/B dadda_fa_4_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/CIN dadda_fa_5_70_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_86_2 U$$2307/X U$$2440/X U$$2573/X VGND VGND VPWR VPWR dadda_fa_2_87_3/B
+ dadda_fa_2_86_5/A sky130_fd_sc_hd__fa_1
XFILLER_131_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_63_1 dadda_fa_4_63_1/A dadda_fa_4_63_1/B dadda_fa_4_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/B dadda_fa_5_63_1/B sky130_fd_sc_hd__fa_1
XFILLER_89_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_79_1 U$$1495/X U$$1628/X U$$1761/X VGND VGND VPWR VPWR dadda_fa_2_80_0/CIN
+ dadda_fa_2_79_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_40_0 dadda_fa_7_40_0/A dadda_fa_7_40_0/B dadda_fa_7_40_0/CIN VGND VGND
+ VPWR VPWR _465_/D _336_/D sky130_fd_sc_hd__fa_1
XFILLER_58_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_56_0 dadda_fa_4_56_0/A dadda_fa_4_56_0/B dadda_fa_4_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/A dadda_fa_5_56_1/A sky130_fd_sc_hd__fa_1
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$210 final_adder.U$$705/A final_adder.U$$704/A VGND VGND VPWR VPWR
+ final_adder.U$$296/A sky130_fd_sc_hd__and2_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$221 final_adder.U$$715/A final_adder.U$$587/B1 final_adder.U$$221/B1
+ VGND VGND VPWR VPWR final_adder.U$$221/X sky130_fd_sc_hd__a21o_1
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$232 final_adder.U$$727/A final_adder.U$$726/A VGND VGND VPWR VPWR
+ final_adder.U$$308/B sky130_fd_sc_hd__and2_1
XFILLER_58_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$243 final_adder.U$$737/A final_adder.U$$609/B1 final_adder.U$$243/B1
+ VGND VGND VPWR VPWR final_adder.U$$243/X sky130_fd_sc_hd__a21o_1
XFILLER_57_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$104 U$$650/B1 U$$118/A2 U$$515/B1 U$$118/B2 VGND VGND VPWR VPWR U$$105/A sky130_fd_sc_hd__a22o_1
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$265 final_adder.U$$264/A final_adder.U$$145/X final_adder.U$$147/X
+ VGND VGND VPWR VPWR final_adder.U$$265/X sky130_fd_sc_hd__a21o_1
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$276 final_adder.U$$276/A final_adder.U$$276/B VGND VGND VPWR VPWR
+ final_adder.U$$330/B sky130_fd_sc_hd__and2_1
Xrepeater480 U$$3537/A2 VGND VGND VPWR VPWR U$$3519/A2 sky130_fd_sc_hd__buf_4
XU$$115 U$$115/A U$$117/B VGND VGND VPWR VPWR U$$115/X sky130_fd_sc_hd__xor2_1
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_530_ _530_/CLK _530_/D VGND VGND VPWR VPWR _530_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$287 final_adder.U$$286/A final_adder.U$$189/X final_adder.U$$191/X
+ VGND VGND VPWR VPWR final_adder.U$$287/X sky130_fd_sc_hd__a21o_1
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$126 U$$811/A1 U$$128/A2 U$$676/A1 U$$128/B2 VGND VGND VPWR VPWR U$$127/A sky130_fd_sc_hd__a22o_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater491 U$$3404/A2 VGND VGND VPWR VPWR U$$3402/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$298 final_adder.U$$298/A final_adder.U$$298/B VGND VGND VPWR VPWR
+ final_adder.U$$340/A sky130_fd_sc_hd__and2_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$137 U$$2/A VGND VGND VPWR VPWR U$$137/Y sky130_fd_sc_hd__inv_1
XFILLER_72_334 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$148 U$$148/A U$$180/B VGND VGND VPWR VPWR U$$148/X sky130_fd_sc_hd__xor2_1
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$159 U$$707/A1 U$$175/A2 U$$22/B1 U$$175/B2 VGND VGND VPWR VPWR U$$160/A sky130_fd_sc_hd__a22o_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_461_ _463_/CLK _461_/D VGND VGND VPWR VPWR _461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_392_ _521_/CLK _392_/D VGND VGND VPWR VPWR _392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1004 _657_/Q VGND VGND VPWR VPWR U$$2861/B sky130_fd_sc_hd__buf_6
Xrepeater1015 U$$2708/B VGND VGND VPWR VPWR U$$2706/B sky130_fd_sc_hd__buf_6
Xrepeater1026 _653_/Q VGND VGND VPWR VPWR U$$2583/B sky130_fd_sc_hd__buf_6
XFILLER_153_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1037 _651_/Q VGND VGND VPWR VPWR U$$2466/A sky130_fd_sc_hd__buf_6
Xrepeater1048 U$$2174/B VGND VGND VPWR VPWR U$$2136/B sky130_fd_sc_hd__buf_6
XFILLER_107_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1059 U$$2039/B VGND VGND VPWR VPWR U$$2029/B sky130_fd_sc_hd__buf_8
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_74_0 dadda_fa_0_74_0/A U$$820/X U$$953/X VGND VGND VPWR VPWR dadda_fa_1_75_7/CIN
+ dadda_fa_1_74_8/B sky130_fd_sc_hd__fa_1
XFILLER_96_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput250 c[94] VGND VGND VPWR VPWR input250/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_194 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$660 U$$934/A1 U$$668/A2 U$$936/A1 U$$670/B2 VGND VGND VPWR VPWR U$$661/A sky130_fd_sc_hd__a22o_1
X_659_ _674_/CLK _659_/D VGND VGND VPWR VPWR _659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$671 U$$671/A U$$685/A VGND VGND VPWR VPWR U$$671/X sky130_fd_sc_hd__xor2_1
XFILLER_56_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$682 U$$817/B1 U$$682/A2 U$$682/B1 U$$682/B2 VGND VGND VPWR VPWR U$$683/A sky130_fd_sc_hd__a22o_1
XU$$693 U$$828/B1 U$$759/A2 U$$695/A1 U$$759/B2 VGND VGND VPWR VPWR U$$694/A sky130_fd_sc_hd__a22o_1
XFILLER_210_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1239_1715 VGND VGND VPWR VPWR U$$1239_1715/HI U$$1239/A1 sky130_fd_sc_hd__conb_1
XFILLER_117_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_80_1 dadda_fa_5_80_1/A dadda_fa_5_80_1/B dadda_fa_5_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_81_0/B dadda_fa_7_80_0/A sky130_fd_sc_hd__fa_2
XFILLER_172_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_96_1 U$$2859/X U$$2992/X U$$3125/X VGND VGND VPWR VPWR dadda_fa_3_97_0/CIN
+ dadda_fa_3_96_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_73_0 dadda_fa_5_73_0/A dadda_fa_5_73_0/B dadda_fa_5_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_74_0/A dadda_fa_6_73_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1560 U$$4291/A1 VGND VGND VPWR VPWR U$$3741/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_89_0 U$$3377/X U$$3510/X U$$3643/X VGND VGND VPWR VPWR dadda_fa_3_90_0/B
+ dadda_fa_3_89_2/B sky130_fd_sc_hd__fa_1
XFILLER_119_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1571 U$$451/A1 VGND VGND VPWR VPWR U$$449/B1 sky130_fd_sc_hd__buf_6
Xrepeater1582 U$$584/B1 VGND VGND VPWR VPWR U$$3187/B1 sky130_fd_sc_hd__buf_6
Xrepeater1593 U$$4418/B1 VGND VGND VPWR VPWR U$$2774/B1 sky130_fd_sc_hd__buf_4
XFILLER_63_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_72_8 dadda_fa_1_72_8/A dadda_fa_1_72_8/B dadda_fa_1_72_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_73_3/A dadda_fa_3_72_0/A sky130_fd_sc_hd__fa_2
XFILLER_101_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_65_7 dadda_fa_1_65_7/A dadda_fa_1_65_7/B dadda_fa_1_65_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_2/CIN dadda_fa_2_65_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_6 U$$3980/X U$$4036/B input210/X VGND VGND VPWR VPWR dadda_fa_2_59_2/B
+ dadda_fa_2_58_5/B sky130_fd_sc_hd__fa_1
XFILLER_66_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_92_2 U$$2718/X U$$2851/X VGND VGND VPWR VPWR dadda_fa_2_93_5/B dadda_fa_3_92_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_88_0 dadda_fa_7_88_0/A dadda_fa_7_88_0/B dadda_fa_7_88_0/CIN VGND VGND
+ VPWR VPWR _513_/D _384_/D sky130_fd_sc_hd__fa_1
XFILLER_136_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_91_0 U$$1917/Y U$$2051/X U$$2184/X VGND VGND VPWR VPWR dadda_fa_2_92_4/B
+ dadda_fa_2_91_5/B sky130_fd_sc_hd__fa_1
XFILLER_11_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4408 U$$4408/A1 U$$4388/X _561_/Q U$$4430/B2 VGND VGND VPWR VPWR U$$4409/A sky130_fd_sc_hd__a22o_1
XU$$4419 U$$4419/A U$$4419/B VGND VGND VPWR VPWR U$$4419/X sky130_fd_sc_hd__xor2_1
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3707 U$$3844/A1 U$$3743/A2 _553_/Q U$$3743/B2 VGND VGND VPWR VPWR U$$3708/A sky130_fd_sc_hd__a22o_1
XFILLER_46_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3718 U$$3718/A U$$3740/B VGND VGND VPWR VPWR U$$3718/X sky130_fd_sc_hd__xor2_1
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3729 U$$4003/A1 U$$3833/A2 _564_/Q U$$3833/B2 VGND VGND VPWR VPWR U$$3730/A sky130_fd_sc_hd__a22o_1
XFILLER_38_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_103_0 dadda_fa_6_103_0/A dadda_fa_6_103_0/B dadda_fa_6_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_104_0/B dadda_fa_7_103_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1778_1724 VGND VGND VPWR VPWR U$$1778_1724/HI U$$1778/B1 sky130_fd_sc_hd__conb_1
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_300 _235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_311 _236_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_322 _238_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_513_ _514_/CLK _513_/D VGND VGND VPWR VPWR _513_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 _239_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_23_3 U$$1516/X input172/X dadda_fa_3_23_3/CIN VGND VGND VPWR VPWR dadda_fa_4_24_1/B
+ dadda_fa_4_23_2/CIN sky130_fd_sc_hd__fa_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_344 U$$80/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_355 U$$3735/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_366 _554_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_444_ _444_/CLK _444_/D VGND VGND VPWR VPWR _444_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_377 U$$811/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_388 _564_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_310 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_375_ _507_/CLK _375_/D VGND VGND VPWR VPWR _375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1070 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_90_0 dadda_fa_6_90_0/A dadda_fa_6_90_0/B dadda_fa_6_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_91_0/B dadda_fa_7_90_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_103_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_68_5 dadda_fa_2_68_5/A dadda_fa_2_68_5/B dadda_fa_2_68_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_2/A dadda_fa_4_68_0/A sky130_fd_sc_hd__fa_1
XFILLER_96_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$490 U$$490/A U$$532/B VGND VGND VPWR VPWR U$$490/X sky130_fd_sc_hd__xor2_1
XFILLER_211_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_623 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1390 U$$4194/B1 VGND VGND VPWR VPWR U$$3783/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_70_5 U$$4270/X U$$4403/X input224/X VGND VGND VPWR VPWR dadda_fa_2_71_2/A
+ dadda_fa_2_70_5/A sky130_fd_sc_hd__fa_1
XFILLER_101_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_63_4 U$$3990/X U$$4123/X U$$4256/X VGND VGND VPWR VPWR dadda_fa_2_64_1/CIN
+ dadda_fa_2_63_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_56_3 U$$2380/X U$$2513/X U$$2646/X VGND VGND VPWR VPWR dadda_fa_2_57_1/B
+ dadda_fa_2_56_4/B sky130_fd_sc_hd__fa_1
XFILLER_132_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_33_2 dadda_fa_4_33_2/A dadda_fa_4_33_2/B dadda_fa_4_33_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/CIN dadda_fa_5_33_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_41_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_49_2 U$$903/X U$$1036/X U$$1169/X VGND VGND VPWR VPWR dadda_fa_2_50_1/B
+ dadda_fa_2_49_4/B sky130_fd_sc_hd__fa_1
XFILLER_54_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_26_1 dadda_fa_4_26_1/A dadda_fa_4_26_1/B dadda_fa_4_26_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/B dadda_fa_5_26_1/B sky130_fd_sc_hd__fa_1
XFILLER_199_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_19_0 U$$1109/X U$$1242/X input167/X VGND VGND VPWR VPWR dadda_fa_5_20_0/A
+ dadda_fa_5_19_1/A sky130_fd_sc_hd__fa_1
XFILLER_199_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4205 U$$4205/A U$$4247/A VGND VGND VPWR VPWR U$$4205/X sky130_fd_sc_hd__xor2_1
XU$$4216 U$$4353/A1 U$$4244/A2 U$$4218/A1 U$$4244/B2 VGND VGND VPWR VPWR U$$4217/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4227 U$$4227/A U$$4239/B VGND VGND VPWR VPWR U$$4227/X sky130_fd_sc_hd__xor2_1
XFILLER_59_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4238 U$$4238/A1 U$$4238/A2 U$$4238/B1 U$$4238/B2 VGND VGND VPWR VPWR U$$4239/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3504 U$$3504/A U$$3506/B VGND VGND VPWR VPWR U$$3504/X sky130_fd_sc_hd__xor2_1
XFILLER_65_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4249 U$$4350/B VGND VGND VPWR VPWR U$$4249/Y sky130_fd_sc_hd__inv_1
XU$$3515 U$$3652/A1 U$$3537/A2 U$$3789/B1 U$$3537/B2 VGND VGND VPWR VPWR U$$3516/A
+ sky130_fd_sc_hd__a22o_1
XU$$3526 U$$3526/A U$$3538/B VGND VGND VPWR VPWR U$$3526/X sky130_fd_sc_hd__xor2_1
XFILLER_74_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3537 _604_/Q U$$3537/A2 U$$3539/A1 U$$3537/B2 VGND VGND VPWR VPWR U$$3538/A sky130_fd_sc_hd__a22o_1
XFILLER_46_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2803 U$$2803/A U$$2839/B VGND VGND VPWR VPWR U$$2803/X sky130_fd_sc_hd__xor2_1
XU$$3548 U$$3548/A U$$3556/B VGND VGND VPWR VPWR U$$3548/X sky130_fd_sc_hd__xor2_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2814 U$$4184/A1 U$$2814/A2 U$$896/B1 U$$2814/B2 VGND VGND VPWR VPWR U$$2815/A
+ sky130_fd_sc_hd__a22o_1
XU$$3559 U$$4105/B1 U$$3559/A2 U$$3559/B1 U$$3559/B2 VGND VGND VPWR VPWR U$$3560/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2825 U$$2825/A U$$2827/B VGND VGND VPWR VPWR U$$2825/X sky130_fd_sc_hd__xor2_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2836 U$$2971/B1 U$$2744/X U$$2838/A1 U$$2745/X VGND VGND VPWR VPWR U$$2837/A sky130_fd_sc_hd__a22o_1
XFILLER_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2847 U$$2847/A U$$2875/B VGND VGND VPWR VPWR U$$2847/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_21_0 U$$49/X U$$182/X U$$315/X VGND VGND VPWR VPWR dadda_fa_4_22_0/B dadda_fa_4_21_1/CIN
+ sky130_fd_sc_hd__fa_1
XANTENNA_130 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2858 U$$2858/A1 U$$2866/A2 _608_/Q U$$2866/B2 VGND VGND VPWR VPWR U$$2859/A sky130_fd_sc_hd__a22o_1
XFILLER_33_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2869 U$$2869/A _657_/Q VGND VGND VPWR VPWR U$$2869/X sky130_fd_sc_hd__xor2_1
XANTENNA_152 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 _183_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_551 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_196 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_427_ _428_/CLK _427_/D VGND VGND VPWR VPWR _427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_358_ _487_/CLK _358_/D VGND VGND VPWR VPWR _358_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_289_ _526_/CLK _289_/D VGND VGND VPWR VPWR _289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_80_4 dadda_fa_2_80_4/A dadda_fa_2_80_4/B dadda_fa_2_80_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/CIN dadda_fa_3_80_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_73_3 dadda_fa_2_73_3/A dadda_fa_2_73_3/B dadda_fa_2_73_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/B dadda_fa_3_73_3/B sky130_fd_sc_hd__fa_1
XFILLER_29_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_66_2 dadda_fa_2_66_2/A dadda_fa_2_66_2/B dadda_fa_2_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/A dadda_fa_3_66_3/A sky130_fd_sc_hd__fa_2
XFILLER_116_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_43_1 dadda_fa_5_43_1/A dadda_fa_5_43_1/B dadda_fa_5_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_44_0/B dadda_fa_7_43_0/A sky130_fd_sc_hd__fa_2
XFILLER_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_59_1 dadda_fa_2_59_1/A dadda_fa_2_59_1/B dadda_fa_2_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_0/CIN dadda_fa_3_59_2/CIN sky130_fd_sc_hd__fa_1
Xinput3 a[11] VGND VGND VPWR VPWR _627_/D sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_5_36_0 dadda_fa_5_36_0/A dadda_fa_5_36_0/B dadda_fa_5_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_37_0/A dadda_fa_6_36_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_37_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4421_1789 VGND VGND VPWR VPWR U$$4421_1789/HI U$$4421/B sky130_fd_sc_hd__conb_1
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_110_0 dadda_fa_5_110_0/A dadda_fa_5_110_0/B dadda_fa_5_110_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_111_0/A dadda_fa_6_110_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_203_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1 _425_/Q _297_/Q VGND VGND VPWR VPWR final_adder.U$$129/B1 final_adder.U$$623/A
+ sky130_fd_sc_hd__ha_1
XFILLER_152_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput340 _173_/Q VGND VGND VPWR VPWR o[5] sky130_fd_sc_hd__buf_2
XFILLER_82_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput351 _174_/Q VGND VGND VPWR VPWR o[6] sky130_fd_sc_hd__buf_2
Xoutput362 _175_/Q VGND VGND VPWR VPWR o[7] sky130_fd_sc_hd__buf_2
XFILLER_160_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput373 _176_/Q VGND VGND VPWR VPWR o[8] sky130_fd_sc_hd__buf_2
XFILLER_156_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput384 _177_/Q VGND VGND VPWR VPWR o[9] sky130_fd_sc_hd__buf_2
XFILLER_102_832 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_61_1 U$$2390/X U$$2523/X U$$2656/X VGND VGND VPWR VPWR dadda_fa_2_62_0/CIN
+ dadda_fa_2_61_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_0 U$$780/X U$$913/X U$$1046/X VGND VGND VPWR VPWR dadda_fa_2_55_0/B
+ dadda_fa_2_54_3/B sky130_fd_sc_hd__fa_1
XFILLER_142_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_941 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1409 U$$1409/A U$$1443/B VGND VGND VPWR VPWR U$$1409/X sky130_fd_sc_hd__xor2_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_212_ _213_/CLK _212_/D VGND VGND VPWR VPWR _212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_90_3 dadda_fa_3_90_3/A dadda_fa_3_90_3/B dadda_fa_3_90_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_1/B dadda_fa_4_90_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_183_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_721 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_83_2 dadda_fa_3_83_2/A dadda_fa_3_83_2/B dadda_fa_3_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_1/A dadda_fa_4_83_2/B sky130_fd_sc_hd__fa_1
XFILLER_87_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_76_1 dadda_fa_3_76_1/A dadda_fa_3_76_1/B dadda_fa_3_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_0/CIN dadda_fa_4_76_2/A sky130_fd_sc_hd__fa_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_53_0 dadda_fa_6_53_0/A dadda_fa_6_53_0/B dadda_fa_6_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_54_0/B dadda_fa_7_53_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_69_0 dadda_fa_3_69_0/A dadda_fa_3_69_0/B dadda_fa_3_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_0/B dadda_fa_4_69_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4002 U$$4002/A U$$4036/B VGND VGND VPWR VPWR U$$4002/X sky130_fd_sc_hd__xor2_1
XU$$4013 U$$4287/A1 U$$4029/A2 _569_/Q U$$4029/B2 VGND VGND VPWR VPWR U$$4014/A sky130_fd_sc_hd__a22o_1
XU$$4024 U$$4024/A U$$4044/B VGND VGND VPWR VPWR U$$4024/X sky130_fd_sc_hd__xor2_1
XFILLER_47_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4035 U$$4035/A1 U$$4035/A2 U$$4035/B1 U$$4081/B2 VGND VGND VPWR VPWR U$$4036/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_700 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3301 U$$3301/A U$$3363/B VGND VGND VPWR VPWR U$$3301/X sky130_fd_sc_hd__xor2_1
XU$$4046 U$$4046/A U$$4070/B VGND VGND VPWR VPWR U$$4046/X sky130_fd_sc_hd__xor2_1
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4057 _590_/Q U$$4061/A2 U$$4194/B1 U$$4061/B2 VGND VGND VPWR VPWR U$$4058/A sky130_fd_sc_hd__a22o_1
XU$$3312 U$$3447/B1 U$$3356/A2 U$$3312/B1 U$$3356/B2 VGND VGND VPWR VPWR U$$3313/A
+ sky130_fd_sc_hd__a22o_1
XU$$4068 U$$4068/A U$$4070/B VGND VGND VPWR VPWR U$$4068/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_2 dadda_fa_4_112_2/A dadda_fa_4_112_2/B dadda_ha_3_112_2/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_113_0/CIN dadda_fa_5_112_1/CIN sky130_fd_sc_hd__fa_1
XU$$3323 U$$3323/A U$$3369/B VGND VGND VPWR VPWR U$$3323/X sky130_fd_sc_hd__xor2_1
XU$$3334 U$$4430/A1 U$$3368/A2 U$$4432/A1 U$$3368/B2 VGND VGND VPWR VPWR U$$3335/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4079 U$$4353/A1 U$$3977/X U$$4218/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4080/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2600 U$$2872/B1 U$$2600/A2 U$$2600/B1 U$$2600/B2 VGND VGND VPWR VPWR U$$2601/A
+ sky130_fd_sc_hd__a22o_1
XU$$3345 U$$3345/A U$$3363/B VGND VGND VPWR VPWR U$$3345/X sky130_fd_sc_hd__xor2_1
XFILLER_46_451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3356 U$$4450/B1 U$$3356/A2 U$$3358/A1 U$$3356/B2 VGND VGND VPWR VPWR U$$3357/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2611 U$$2611/A1 U$$2697/A2 U$$2611/B1 U$$2697/B2 VGND VGND VPWR VPWR U$$2612/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2622 U$$2622/A U$$2654/B VGND VGND VPWR VPWR U$$2622/X sky130_fd_sc_hd__xor2_1
XU$$3367 U$$3367/A U$$3424/A VGND VGND VPWR VPWR U$$3367/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_105_1 dadda_fa_4_105_1/A dadda_fa_4_105_1/B dadda_fa_4_105_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/B dadda_fa_5_105_1/B sky130_fd_sc_hd__fa_1
XFILLER_111_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2633 U$$715/A1 U$$2687/A2 U$$3181/B1 U$$2687/B2 VGND VGND VPWR VPWR U$$2634/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3378 U$$4198/B1 U$$3378/A2 U$$3380/A1 U$$3378/B2 VGND VGND VPWR VPWR U$$3379/A
+ sky130_fd_sc_hd__a22o_1
XU$$2644 U$$2644/A U$$2688/B VGND VGND VPWR VPWR U$$2644/X sky130_fd_sc_hd__xor2_1
XFILLER_206_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3389 U$$3389/A U$$3397/B VGND VGND VPWR VPWR U$$3389/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1910 U$$1910/A U$$1918/A VGND VGND VPWR VPWR U$$1910/X sky130_fd_sc_hd__xor2_1
XFILLER_62_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2655 U$$463/A1 U$$2663/A2 U$$54/A1 U$$2663/B2 VGND VGND VPWR VPWR U$$2656/A sky130_fd_sc_hd__a22o_1
XU$$2666 U$$2666/A U$$2706/B VGND VGND VPWR VPWR U$$2666/X sky130_fd_sc_hd__xor2_1
XU$$1921 _645_/Q U$$1921/B VGND VGND VPWR VPWR U$$1921/X sky130_fd_sc_hd__and2_1
XFILLER_179_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1932 U$$2343/A1 U$$2010/A2 U$$2345/A1 U$$2010/B2 VGND VGND VPWR VPWR U$$1933/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2677 U$$3362/A1 U$$2697/A2 U$$3362/B1 U$$2697/B2 VGND VGND VPWR VPWR U$$2678/A
+ sky130_fd_sc_hd__a22o_1
XU$$2688 U$$2688/A U$$2688/B VGND VGND VPWR VPWR U$$2688/X sky130_fd_sc_hd__xor2_1
XU$$1943 U$$1943/A U$$1983/B VGND VGND VPWR VPWR U$$1943/X sky130_fd_sc_hd__xor2_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1954 U$$36/A1 U$$1956/A2 U$$997/A1 U$$1956/B2 VGND VGND VPWR VPWR U$$1955/A sky130_fd_sc_hd__a22o_1
XFILLER_62_999 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2699 U$$3245/B1 U$$2707/A2 U$$3112/A1 U$$2707/B2 VGND VGND VPWR VPWR U$$2700/A
+ sky130_fd_sc_hd__a22o_1
XU$$1965 U$$1965/A U$$1983/B VGND VGND VPWR VPWR U$$1965/X sky130_fd_sc_hd__xor2_1
XFILLER_15_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1976 U$$1976/A1 U$$1976/A2 U$$3485/A1 U$$1976/B2 VGND VGND VPWR VPWR U$$1977/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_126_0 dadda_fa_7_126_0/A dadda_fa_7_126_0/B dadda_fa_7_126_0/CIN VGND
+ VGND VPWR VPWR _551_/D _422_/D sky130_fd_sc_hd__fa_1
XU$$1987 U$$1987/A U$$2011/B VGND VGND VPWR VPWR U$$1987/X sky130_fd_sc_hd__xor2_1
XFILLER_30_830 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1998 U$$3642/A1 U$$1922/X U$$3505/B1 U$$1923/X VGND VGND VPWR VPWR U$$1999/A sky130_fd_sc_hd__a22o_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_71_0 dadda_fa_2_71_0/A dadda_fa_2_71_0/B dadda_fa_2_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_0/B dadda_fa_3_71_2/B sky130_fd_sc_hd__fa_1
XFILLER_97_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater810 U$$2302/B2 VGND VGND VPWR VPWR U$$2298/B2 sky130_fd_sc_hd__buf_6
Xrepeater821 U$$2185/B2 VGND VGND VPWR VPWR U$$2189/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$617 final_adder.U$$744/A final_adder.U$$744/B final_adder.U$$617/B1
+ VGND VGND VPWR VPWR final_adder.U$$745/B sky130_fd_sc_hd__a21o_1
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$628 final_adder.U$$628/A final_adder.U$$628/B VGND VGND VPWR VPWR
+ _174_/D sky130_fd_sc_hd__xor2_1
Xrepeater832 U$$1851/B2 VGND VGND VPWR VPWR U$$1843/B2 sky130_fd_sc_hd__buf_6
XFILLER_96_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater843 U$$1768/B2 VGND VGND VPWR VPWR U$$1762/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$639 final_adder.U$$639/A final_adder.U$$639/B VGND VGND VPWR VPWR
+ _185_/D sky130_fd_sc_hd__xor2_4
XFILLER_110_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater854 U$$1512/X VGND VGND VPWR VPWR U$$1635/B2 sky130_fd_sc_hd__clkbuf_8
Xrepeater865 U$$1474/B2 VGND VGND VPWR VPWR U$$1458/B2 sky130_fd_sc_hd__buf_4
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater876 U$$1238/X VGND VGND VPWR VPWR U$$1323/B2 sky130_fd_sc_hd__buf_4
Xrepeater887 U$$1101/X VGND VGND VPWR VPWR U$$1208/B2 sky130_fd_sc_hd__buf_6
Xrepeater898 U$$4480/B2 VGND VGND VPWR VPWR U$$4454/B2 sky130_fd_sc_hd__buf_6
XU$$50 U$$50/A1 U$$52/A2 U$$52/A1 U$$52/B2 VGND VGND VPWR VPWR U$$51/A sky130_fd_sc_hd__a22o_1
XU$$61 U$$61/A U$$3/A VGND VGND VPWR VPWR U$$61/X sky130_fd_sc_hd__xor2_1
XFILLER_53_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$72 U$$72/A1 U$$84/A2 U$$74/A1 U$$84/B2 VGND VGND VPWR VPWR U$$73/A sky130_fd_sc_hd__a22o_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$83 U$$83/A U$$85/B VGND VGND VPWR VPWR U$$83/X sky130_fd_sc_hd__xor2_1
XU$$94 U$$94/A1 U$$98/A2 U$$96/A1 U$$98/B2 VGND VGND VPWR VPWR U$$95/A sky130_fd_sc_hd__a22o_1
XU$$3890 U$$4027/A1 U$$3916/A2 _576_/Q U$$3916/B2 VGND VGND VPWR VPWR U$$3891/A sky130_fd_sc_hd__a22o_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_30 _282_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_41 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_835 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_52 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_96 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_93_1 dadda_fa_4_93_1/A dadda_fa_4_93_1/B dadda_fa_4_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/B dadda_fa_5_93_1/B sky130_fd_sc_hd__fa_1
XFILLER_10_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_70_0 dadda_fa_7_70_0/A dadda_fa_7_70_0/B dadda_fa_7_70_0/CIN VGND VGND
+ VPWR VPWR _495_/D _366_/D sky130_fd_sc_hd__fa_1
XFILLER_192_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_86_0 dadda_fa_4_86_0/A dadda_fa_4_86_0/B dadda_fa_4_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/A dadda_fa_5_86_1/A sky130_fd_sc_hd__fa_1
XFILLER_180_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_107_3 input137/X dadda_fa_3_107_3/B dadda_fa_3_107_3/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_108_1/B dadda_fa_4_107_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1206 U$$4357/A1 U$$1208/A2 U$$658/B1 U$$1208/B2 VGND VGND VPWR VPWR U$$1207/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1217 U$$1217/A U$$1232/A VGND VGND VPWR VPWR U$$1217/X sky130_fd_sc_hd__xor2_1
XFILLER_203_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1228 U$$954/A1 U$$1230/A2 U$$817/B1 U$$1230/B2 VGND VGND VPWR VPWR U$$1229/A sky130_fd_sc_hd__a22o_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1239 U$$1239/A1 U$$1323/A2 U$$967/A1 U$$1323/B2 VGND VGND VPWR VPWR U$$1240/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_25 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_50_5 dadda_fa_2_50_5/A dadda_fa_2_50_5/B dadda_fa_2_50_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_2/A dadda_fa_4_50_0/A sky130_fd_sc_hd__fa_1
XFILLER_93_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_43_4 dadda_fa_2_43_4/A dadda_fa_2_43_4/B dadda_fa_2_43_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_1/CIN dadda_fa_3_43_3/CIN sky130_fd_sc_hd__fa_1
XU$$3120 U$$3255/B1 U$$3120/A2 _602_/Q U$$3120/B2 VGND VGND VPWR VPWR U$$3121/A sky130_fd_sc_hd__a22o_1
XFILLER_81_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3131 U$$3131/A U$$3133/B VGND VGND VPWR VPWR U$$3131/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_6_2_0 U$$11/X U$$144/X VGND VGND VPWR VPWR dadda_fa_7_3_0/B dadda_ha_6_2_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$3142 U$$3551/B1 U$$3144/A2 U$$3281/A1 U$$3144/B2 VGND VGND VPWR VPWR U$$3143/A
+ sky130_fd_sc_hd__a22o_1
XU$$3153 U$$3288/A VGND VGND VPWR VPWR U$$3153/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_2_36_3 U$$1941/X U$$2074/X U$$2207/X VGND VGND VPWR VPWR dadda_fa_3_37_1/B
+ dadda_fa_3_36_3/B sky130_fd_sc_hd__fa_1
XFILLER_19_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1504_1720 VGND VGND VPWR VPWR U$$1504_1720/HI U$$1504/B1 sky130_fd_sc_hd__conb_1
XU$$3164 U$$3164/A U$$3232/B VGND VGND VPWR VPWR U$$3164/X sky130_fd_sc_hd__xor2_1
XFILLER_19_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3175 U$$3175/A1 U$$3215/A2 U$$4410/A1 U$$3215/B2 VGND VGND VPWR VPWR U$$3176/A
+ sky130_fd_sc_hd__a22o_1
XU$$2430 U$$2430/A U$$2465/A VGND VGND VPWR VPWR U$$2430/X sky130_fd_sc_hd__xor2_1
XU$$2441 U$$4494/B1 U$$2451/A2 U$$4224/A1 U$$2451/B2 VGND VGND VPWR VPWR U$$2442/A
+ sky130_fd_sc_hd__a22o_1
XU$$3186 U$$3186/A U$$3208/B VGND VGND VPWR VPWR U$$3186/X sky130_fd_sc_hd__xor2_1
XU$$2452 U$$2452/A U$$2465/A VGND VGND VPWR VPWR U$$2452/X sky130_fd_sc_hd__xor2_1
XU$$3197 U$$4430/A1 U$$3235/A2 U$$4432/A1 U$$3235/B2 VGND VGND VPWR VPWR U$$3198/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2463 _615_/Q U$$2463/A2 U$$2463/B1 U$$2463/B2 VGND VGND VPWR VPWR U$$2464/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_29_2 U$$863/X U$$996/X U$$1129/X VGND VGND VPWR VPWR dadda_fa_3_30_2/A
+ dadda_fa_3_29_3/CIN sky130_fd_sc_hd__fa_2
XU$$2474 U$$2611/A1 U$$2516/A2 U$$2611/B1 U$$2516/B2 VGND VGND VPWR VPWR U$$2475/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2485 U$$2485/A U$$2531/B VGND VGND VPWR VPWR U$$2485/X sky130_fd_sc_hd__xor2_1
XU$$1740 U$$3245/B1 U$$1740/A2 U$$3112/A1 U$$1740/B2 VGND VGND VPWR VPWR U$$1741/A
+ sky130_fd_sc_hd__a22o_1
XU$$1751 U$$1751/A U$$1763/B VGND VGND VPWR VPWR U$$1751/X sky130_fd_sc_hd__xor2_1
XU$$2496 U$$4140/A1 U$$2516/A2 U$$3181/B1 U$$2516/B2 VGND VGND VPWR VPWR U$$2497/A
+ sky130_fd_sc_hd__a22o_1
XU$$1762 U$$253/B1 U$$1762/A2 U$$2721/B1 U$$1762/B2 VGND VGND VPWR VPWR U$$1763/A
+ sky130_fd_sc_hd__a22o_1
XU$$1773 U$$1773/A U$$1773/B VGND VGND VPWR VPWR U$$1773/X sky130_fd_sc_hd__xor2_1
XU$$1784 U$$1918/A U$$1784/B VGND VGND VPWR VPWR U$$1784/X sky130_fd_sc_hd__and2_1
XFILLER_166_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1795 U$$973/A1 U$$1859/A2 U$$838/A1 U$$1859/B2 VGND VGND VPWR VPWR U$$1796/A sky130_fd_sc_hd__a22o_1
XFILLER_188_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput50 a[54] VGND VGND VPWR VPWR _670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_190_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput61 a[6] VGND VGND VPWR VPWR _622_/D sky130_fd_sc_hd__clkbuf_2
Xinput72 b[16] VGND VGND VPWR VPWR _568_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_721 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput83 b[26] VGND VGND VPWR VPWR _578_/D sky130_fd_sc_hd__clkbuf_1
Xinput94 b[36] VGND VGND VPWR VPWR _588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1069 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$403 final_adder.U$$348/X final_adder.U$$734/B final_adder.U$$349/X
+ VGND VGND VPWR VPWR final_adder.U$$742/B sky130_fd_sc_hd__a21o_2
XFILLER_85_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$425 final_adder.U$$342/B final_adder.U$$710/B final_adder.U$$301/X
+ VGND VGND VPWR VPWR final_adder.U$$714/B sky130_fd_sc_hd__a21o_1
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater640 U$$1065/B2 VGND VGND VPWR VPWR U$$995/B2 sky130_fd_sc_hd__buf_4
XFILLER_111_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$447 final_adder.U$$270/B final_adder.U$$650/B final_adder.U$$157/X
+ VGND VGND VPWR VPWR final_adder.U$$652/B sky130_fd_sc_hd__a21o_1
Xrepeater651 U$$896/B2 VGND VGND VPWR VPWR U$$906/B2 sky130_fd_sc_hd__buf_4
XFILLER_123_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater662 U$$690/X VGND VGND VPWR VPWR U$$795/B2 sky130_fd_sc_hd__buf_4
XFILLER_45_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$469 final_adder.U$$292/B final_adder.U$$694/B final_adder.U$$201/X
+ VGND VGND VPWR VPWR final_adder.U$$696/B sky130_fd_sc_hd__a21o_1
XU$$308 U$$34/A1 U$$308/A2 U$$856/B1 U$$308/B2 VGND VGND VPWR VPWR U$$309/A sky130_fd_sc_hd__a22o_1
XFILLER_85_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater673 U$$4345/B2 VGND VGND VPWR VPWR U$$4297/B2 sky130_fd_sc_hd__buf_6
XFILLER_123_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater684 U$$416/X VGND VGND VPWR VPWR U$$491/B2 sky130_fd_sc_hd__buf_4
XFILLER_38_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$319 U$$319/A U$$319/B VGND VGND VPWR VPWR U$$319/X sky130_fd_sc_hd__xor2_1
XFILLER_38_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater695 U$$4081/B2 VGND VGND VPWR VPWR U$$4005/B2 sky130_fd_sc_hd__buf_4
XFILLER_199_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_914 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_334 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_315 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1208 U$$950/B1 VGND VGND VPWR VPWR U$$676/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_3_112_1 U$$3689/X U$$3822/X U$$3955/X VGND VGND VPWR VPWR dadda_fa_4_113_1/CIN
+ dadda_fa_4_112_2/B sky130_fd_sc_hd__fa_1
Xrepeater1219 U$$4512/A1 VGND VGND VPWR VPWR U$$4238/A1 sky130_fd_sc_hd__buf_6
XFILLER_113_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_105_0 U$$3675/X U$$3808/X U$$3941/X VGND VGND VPWR VPWR dadda_fa_4_106_0/B
+ dadda_fa_4_105_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_53_3 dadda_fa_3_53_3/A dadda_fa_3_53_3/B dadda_fa_3_53_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_1/B dadda_fa_4_53_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_69_3 U$$1608/X U$$1741/X U$$1874/X VGND VGND VPWR VPWR dadda_fa_1_70_7/A
+ dadda_fa_1_69_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_46_2 dadda_fa_3_46_2/A dadda_fa_3_46_2/B dadda_fa_3_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_1/A dadda_fa_4_46_2/B sky130_fd_sc_hd__fa_1
XTAP_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$820 U$$820/A U$$821/A VGND VGND VPWR VPWR U$$820/X sky130_fd_sc_hd__xor2_1
XFILLER_1_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_675_ _679_/CLK _675_/D VGND VGND VPWR VPWR _675_/Q sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_3_39_1 dadda_fa_3_39_1/A dadda_fa_3_39_1/B dadda_fa_3_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_0/CIN dadda_fa_4_39_2/A sky130_fd_sc_hd__fa_1
XU$$831 U$$831/A U$$859/B VGND VGND VPWR VPWR U$$831/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$842 U$$20/A1 U$$878/A2 U$$22/A1 U$$878/B2 VGND VGND VPWR VPWR U$$843/A sky130_fd_sc_hd__a22o_1
XFILLER_204_500 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_16_0 dadda_fa_6_16_0/A dadda_fa_6_16_0/B dadda_fa_6_16_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_17_0/B dadda_fa_7_16_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_44_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$853 U$$853/A U$$925/B VGND VGND VPWR VPWR U$$853/X sky130_fd_sc_hd__xor2_1
XFILLER_90_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1003 U$$2508/B1 U$$979/A2 U$$2375/A1 U$$979/B2 VGND VGND VPWR VPWR U$$1004/A sky130_fd_sc_hd__a22o_1
XFILLER_21_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$864 U$$999/B1 U$$924/A2 U$$866/A1 U$$924/B2 VGND VGND VPWR VPWR U$$865/A sky130_fd_sc_hd__a22o_1
XFILLER_56_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$875 U$$875/A U$$879/B VGND VGND VPWR VPWR U$$875/X sky130_fd_sc_hd__xor2_1
XU$$1014 U$$1014/A U$$982/B VGND VGND VPWR VPWR U$$1014/X sky130_fd_sc_hd__xor2_1
XU$$886 U$$64/A1 U$$928/A2 U$$66/A1 U$$928/B2 VGND VGND VPWR VPWR U$$887/A sky130_fd_sc_hd__a22o_1
XU$$1025 U$$749/B1 U$$997/A2 U$$68/A1 U$$997/B2 VGND VGND VPWR VPWR U$$1026/A sky130_fd_sc_hd__a22o_1
XFILLER_95_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1036 U$$1036/A U$$1040/B VGND VGND VPWR VPWR U$$1036/X sky130_fd_sc_hd__xor2_1
XFILLER_32_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$897 U$$897/A U$$897/B VGND VGND VPWR VPWR U$$897/X sky130_fd_sc_hd__xor2_1
XU$$1047 U$$910/A1 U$$1089/A2 U$$912/A1 U$$1089/B2 VGND VGND VPWR VPWR U$$1048/A sky130_fd_sc_hd__a22o_1
XU$$1058 U$$1058/A U$$998/B VGND VGND VPWR VPWR U$$1058/X sky130_fd_sc_hd__xor2_1
XFILLER_73_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1069 U$$932/A1 U$$963/X U$$934/A1 U$$964/X VGND VGND VPWR VPWR U$$1070/A sky130_fd_sc_hd__a22o_1
XFILLER_148_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1020 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_41_1 U$$1951/X U$$2084/X U$$2217/X VGND VGND VPWR VPWR dadda_fa_3_42_0/CIN
+ dadda_fa_3_41_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_34_0 U$$341/X U$$474/X U$$607/X VGND VGND VPWR VPWR dadda_fa_3_35_0/B
+ dadda_fa_3_34_2/B sky130_fd_sc_hd__fa_1
XFILLER_19_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2260 U$$66/B1 U$$2262/A2 U$$890/B1 U$$2262/B2 VGND VGND VPWR VPWR U$$2261/A sky130_fd_sc_hd__a22o_1
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2271 U$$2271/A U$$2309/B VGND VGND VPWR VPWR U$$2271/X sky130_fd_sc_hd__xor2_1
XU$$2282 U$$2830/A1 U$$2298/A2 U$$914/A1 U$$2298/B2 VGND VGND VPWR VPWR U$$2283/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2293 U$$2293/A U$$2321/B VGND VGND VPWR VPWR U$$2293/X sky130_fd_sc_hd__xor2_1
XFILLER_195_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1570 U$$1570/A U$$1578/B VGND VGND VPWR VPWR U$$1570/X sky130_fd_sc_hd__xor2_1
XFILLER_22_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1581 U$$4184/A1 U$$1627/A2 U$$896/B1 U$$1627/B2 VGND VGND VPWR VPWR U$$1582/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1592 U$$1592/A U$$1598/B VGND VGND VPWR VPWR U$$1592/X sky130_fd_sc_hd__xor2_1
XFILLER_50_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_86_3 U$$2706/X U$$2839/X U$$2972/X VGND VGND VPWR VPWR dadda_fa_2_87_3/CIN
+ dadda_fa_2_86_5/B sky130_fd_sc_hd__fa_1
XFILLER_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_63_2 dadda_fa_4_63_2/A dadda_fa_4_63_2/B dadda_fa_4_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/CIN dadda_fa_5_63_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_79_2 U$$1894/X U$$2027/X U$$2160/X VGND VGND VPWR VPWR dadda_fa_2_80_1/A
+ dadda_fa_2_79_4/A sky130_fd_sc_hd__fa_1
XFILLER_103_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_56_1 dadda_fa_4_56_1/A dadda_fa_4_56_1/B dadda_fa_4_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/B dadda_fa_5_56_1/B sky130_fd_sc_hd__fa_1
XFILLER_103_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$200 final_adder.U$$695/A final_adder.U$$694/A VGND VGND VPWR VPWR
+ final_adder.U$$292/B sky130_fd_sc_hd__and2_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$211 final_adder.U$$705/A final_adder.U$$577/B1 final_adder.U$$211/B1
+ VGND VGND VPWR VPWR final_adder.U$$211/X sky130_fd_sc_hd__a21o_1
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_33_0 dadda_fa_7_33_0/A dadda_fa_7_33_0/B dadda_fa_7_33_0/CIN VGND VGND
+ VPWR VPWR _458_/D _329_/D sky130_fd_sc_hd__fa_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk _634_/CLK VGND VGND VPWR VPWR _623_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_97_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$222 final_adder.U$$717/A final_adder.U$$716/A VGND VGND VPWR VPWR
+ final_adder.U$$302/A sky130_fd_sc_hd__and2_1
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_49_0 dadda_fa_4_49_0/A dadda_fa_4_49_0/B dadda_fa_4_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/A dadda_fa_5_49_1/A sky130_fd_sc_hd__fa_1
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$233 final_adder.U$$727/A final_adder.U$$599/B1 final_adder.U$$233/B1
+ VGND VGND VPWR VPWR final_adder.U$$233/X sky130_fd_sc_hd__a21o_1
XFILLER_44_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$244 final_adder.U$$739/A final_adder.U$$738/A VGND VGND VPWR VPWR
+ final_adder.U$$314/B sky130_fd_sc_hd__and2_1
XFILLER_45_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_899 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$105 U$$105/A U$$117/B VGND VGND VPWR VPWR U$$105/X sky130_fd_sc_hd__xor2_1
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater470 U$$3628/A2 VGND VGND VPWR VPWR U$$3612/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$266 final_adder.U$$266/A final_adder.U$$266/B VGND VGND VPWR VPWR
+ final_adder.U$$324/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$277 final_adder.U$$276/A final_adder.U$$169/X final_adder.U$$171/X
+ VGND VGND VPWR VPWR final_adder.U$$277/X sky130_fd_sc_hd__a21o_1
XU$$116 U$$251/B1 U$$118/A2 U$$253/B1 U$$118/B2 VGND VGND VPWR VPWR U$$117/A sky130_fd_sc_hd__a22o_1
Xrepeater481 U$$3537/A2 VGND VGND VPWR VPWR U$$3531/A2 sky130_fd_sc_hd__buf_4
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$127 U$$127/A U$$129/B VGND VGND VPWR VPWR U$$127/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$288 final_adder.U$$288/A final_adder.U$$288/B VGND VGND VPWR VPWR
+ final_adder.U$$336/B sky130_fd_sc_hd__and2_1
XFILLER_79_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater492 U$$3408/A2 VGND VGND VPWR VPWR U$$3404/A2 sky130_fd_sc_hd__buf_6
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$299 final_adder.U$$298/A final_adder.U$$213/X final_adder.U$$215/X
+ VGND VGND VPWR VPWR final_adder.U$$299/X sky130_fd_sc_hd__a21o_1
XU$$138 _618_/Q VGND VGND VPWR VPWR U$$140/B sky130_fd_sc_hd__inv_1
XU$$149 U$$12/A1 U$$181/A2 U$$14/A1 U$$181/B2 VGND VGND VPWR VPWR U$$150/A sky130_fd_sc_hd__a22o_1
XFILLER_72_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_460_ _463_/CLK _460_/D VGND VGND VPWR VPWR _460_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_391_ _519_/CLK _391_/D VGND VGND VPWR VPWR _391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk _432_/CLK VGND VGND VPWR VPWR _466_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1005 U$$2839/B VGND VGND VPWR VPWR U$$2795/B sky130_fd_sc_hd__buf_6
Xrepeater1016 U$$2730/B VGND VGND VPWR VPWR U$$2688/B sky130_fd_sc_hd__buf_6
XFILLER_182_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1027 U$$2603/A VGND VGND VPWR VPWR U$$2597/B sky130_fd_sc_hd__buf_6
XFILLER_4_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1038 U$$2269/B VGND VGND VPWR VPWR U$$2263/B sky130_fd_sc_hd__buf_8
XFILLER_182_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1049 U$$2110/B VGND VGND VPWR VPWR U$$2108/B sky130_fd_sc_hd__buf_8
XFILLER_141_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_74_1 U$$1086/X U$$1219/X U$$1352/X VGND VGND VPWR VPWR dadda_fa_1_75_8/A
+ dadda_fa_1_74_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_51_0 dadda_fa_3_51_0/A dadda_fa_3_51_0/B dadda_fa_3_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_0/B dadda_fa_4_51_1/CIN sky130_fd_sc_hd__fa_1
Xinput240 c[85] VGND VGND VPWR VPWR input240/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_87_clk _628_/CLK VGND VGND VPWR VPWR _547_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput251 c[95] VGND VGND VPWR VPWR input251/X sky130_fd_sc_hd__buf_4
Xdadda_fa_0_67_0 U$$136/Y U$$273/Y U$$407/X VGND VGND VPWR VPWR dadda_fa_1_68_5/B
+ dadda_fa_1_67_7/B sky130_fd_sc_hd__fa_1
XFILLER_49_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_663 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$650 U$$785/B1 U$$650/A2 U$$650/B1 U$$650/B2 VGND VGND VPWR VPWR U$$651/A sky130_fd_sc_hd__a22o_1
X_658_ _660_/CLK _658_/D VGND VGND VPWR VPWR _658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$661 U$$661/A U$$669/B VGND VGND VPWR VPWR U$$661/X sky130_fd_sc_hd__xor2_1
XU$$672 U$$944/B1 U$$552/X U$$674/A1 U$$553/X VGND VGND VPWR VPWR U$$673/A sky130_fd_sc_hd__a22o_1
XU$$683 U$$683/A U$$684/A VGND VGND VPWR VPWR U$$683/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$694 U$$694/A U$$760/B VGND VGND VPWR VPWR U$$694/X sky130_fd_sc_hd__xor2_1
X_589_ _596_/CLK _589_/D VGND VGND VPWR VPWR _589_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_204_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1027 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk _616_/CLK VGND VGND VPWR VPWR _471_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_191_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_96_2 U$$3258/X U$$3391/X U$$3524/X VGND VGND VPWR VPWR dadda_fa_3_97_1/A
+ dadda_fa_3_96_3/A sky130_fd_sc_hd__fa_1
XFILLER_99_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1550 U$$866/B1 VGND VGND VPWR VPWR U$$731/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_73_1 dadda_fa_5_73_1/A dadda_fa_5_73_1/B dadda_fa_5_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_74_0/B dadda_fa_7_73_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_89_1 U$$3776/X U$$3909/X U$$4042/X VGND VGND VPWR VPWR dadda_fa_3_90_0/CIN
+ dadda_fa_3_89_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater1561 _570_/Q VGND VGND VPWR VPWR U$$4291/A1 sky130_fd_sc_hd__buf_8
Xrepeater1572 U$$3054/A1 VGND VGND VPWR VPWR U$$40/A1 sky130_fd_sc_hd__buf_4
Xrepeater1583 _567_/Q VGND VGND VPWR VPWR U$$584/B1 sky130_fd_sc_hd__buf_6
XFILLER_98_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_66_0 dadda_fa_5_66_0/A dadda_fa_5_66_0/B dadda_fa_5_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_67_0/A dadda_fa_6_66_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1594 _566_/Q VGND VGND VPWR VPWR U$$4418/B1 sky130_fd_sc_hd__buf_6
XFILLER_28_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_65_8 dadda_fa_1_65_8/A dadda_fa_1_65_8/B dadda_fa_1_65_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_3/A dadda_fa_3_65_0/A sky130_fd_sc_hd__fa_2
XFILLER_39_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_78_clk _628_/CLK VGND VGND VPWR VPWR _662_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_7 dadda_fa_1_58_7/A dadda_fa_1_58_7/B dadda_fa_1_58_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_59_2/CIN dadda_fa_2_58_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_5_0 U$$283/X input212/X dadda_fa_6_5_0/CIN VGND VGND VPWR VPWR dadda_fa_7_6_0/B
+ dadda_fa_7_5_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2090 U$$2090/A U$$2130/B VGND VGND VPWR VPWR U$$2090/X sky130_fd_sc_hd__xor2_1
XFILLER_211_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_91_1 U$$2317/X U$$2450/X U$$2583/X VGND VGND VPWR VPWR dadda_fa_2_92_4/CIN
+ dadda_fa_2_91_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_85_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_84_0 dadda_fa_1_84_0/A U$$1505/X U$$1638/X VGND VGND VPWR VPWR dadda_fa_2_85_2/A
+ dadda_fa_2_84_4/A sky130_fd_sc_hd__fa_1
XFILLER_46_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$417_1764 VGND VGND VPWR VPWR U$$417_1764/HI U$$417/A1 sky130_fd_sc_hd__conb_1
XFILLER_131_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_69_clk _369_/CLK VGND VGND VPWR VPWR _572_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$4409 U$$4409/A U$$4409/B VGND VGND VPWR VPWR U$$4409/X sky130_fd_sc_hd__xor2_1
XFILLER_161_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_663 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3708 U$$3708/A U$$3760/B VGND VGND VPWR VPWR U$$3708/X sky130_fd_sc_hd__xor2_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3719 U$$4402/B1 U$$3769/A2 U$$4269/A1 U$$3769/B2 VGND VGND VPWR VPWR U$$3720/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1046 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_301 _235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_512_ _560_/CLK _512_/D VGND VGND VPWR VPWR _512_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_312 _236_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_323 _238_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_334 _239_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_345 U$$3096/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_356 _645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_443_ _443_/CLK _443_/D VGND VGND VPWR VPWR _443_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_367 _555_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_378 U$$938/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_389 _565_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_374_ _503_/CLK _374_/D VGND VGND VPWR VPWR _374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_777 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_950 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_83_0 dadda_fa_6_83_0/A dadda_fa_6_83_0/B dadda_fa_6_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_84_0/B dadda_fa_7_83_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_99_0 U$$4461/X input255/X dadda_fa_3_99_0/CIN VGND VGND VPWR VPWR dadda_fa_4_100_0/B
+ dadda_fa_4_99_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_127_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1099 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1004 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$480 U$$480/A U$$484/B VGND VGND VPWR VPWR U$$480/X sky130_fd_sc_hd__xor2_1
XFILLER_211_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$491 U$$491/A1 U$$491/A2 U$$493/A1 U$$491/B2 VGND VGND VPWR VPWR U$$492/A sky130_fd_sc_hd__a22o_1
XFILLER_177_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1102_1713 VGND VGND VPWR VPWR U$$1102_1713/HI U$$1102/A1 sky130_fd_sc_hd__conb_1
XFILLER_146_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1380 U$$3650/A1 VGND VGND VPWR VPWR U$$634/B1 sky130_fd_sc_hd__buf_6
Xrepeater1391 U$$3374/A1 VGND VGND VPWR VPWR U$$86/A1 sky130_fd_sc_hd__buf_4
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_70_6 dadda_fa_1_70_6/A dadda_fa_1_70_6/B dadda_fa_1_70_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_2/B dadda_fa_2_70_5/B sky130_fd_sc_hd__fa_1
XFILLER_140_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_63_5 input216/X dadda_fa_1_63_5/B dadda_fa_1_63_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_64_2/A dadda_fa_2_63_5/A sky130_fd_sc_hd__fa_1
XFILLER_68_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_56_4 U$$2779/X U$$2912/X U$$3045/X VGND VGND VPWR VPWR dadda_fa_2_57_1/CIN
+ dadda_fa_2_56_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_41_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_49_3 U$$1302/X U$$1435/X U$$1568/X VGND VGND VPWR VPWR dadda_fa_2_50_1/CIN
+ dadda_fa_2_49_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_26_2 dadda_fa_4_26_2/A dadda_fa_4_26_2/B dadda_fa_4_26_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/CIN dadda_fa_5_26_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_1 dadda_fa_4_19_1/A dadda_fa_4_19_1/B dadda_fa_4_19_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_20_0/B dadda_fa_5_19_1/B sky130_fd_sc_hd__fa_2
XFILLER_39_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4206 U$$4480/A1 U$$4114/X U$$4206/B1 U$$4115/X VGND VGND VPWR VPWR U$$4207/A sky130_fd_sc_hd__a22o_1
XU$$4217 U$$4217/A U$$4246/A VGND VGND VPWR VPWR U$$4217/X sky130_fd_sc_hd__xor2_1
XFILLER_77_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4228 U$$4500/B1 U$$4238/A2 U$$4228/B1 U$$4238/B2 VGND VGND VPWR VPWR U$$4229/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4239 U$$4239/A U$$4239/B VGND VGND VPWR VPWR U$$4239/X sky130_fd_sc_hd__xor2_1
XU$$3505 U$$3642/A1 U$$3545/A2 U$$3505/B1 U$$3545/B2 VGND VGND VPWR VPWR U$$3506/A
+ sky130_fd_sc_hd__a22o_1
XU$$3516 U$$3516/A U$$3520/B VGND VGND VPWR VPWR U$$3516/X sky130_fd_sc_hd__xor2_1
XFILLER_86_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3527 _599_/Q U$$3531/A2 _600_/Q U$$3531/B2 VGND VGND VPWR VPWR U$$3528/A sky130_fd_sc_hd__a22o_1
XU$$1641_1722 VGND VGND VPWR VPWR U$$1641_1722/HI U$$1641/B1 sky130_fd_sc_hd__conb_1
XFILLER_58_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3538 U$$3538/A U$$3538/B VGND VGND VPWR VPWR U$$3538/X sky130_fd_sc_hd__xor2_1
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3549 U$$4369/B1 U$$3559/A2 U$$4236/A1 U$$3559/B2 VGND VGND VPWR VPWR U$$3550/A
+ sky130_fd_sc_hd__a22o_1
XU$$2804 U$$4035/B1 U$$2832/A2 U$$3902/A1 U$$2832/B2 VGND VGND VPWR VPWR U$$2805/A
+ sky130_fd_sc_hd__a22o_1
XU$$2815 U$$2815/A U$$2827/B VGND VGND VPWR VPWR U$$2815/X sky130_fd_sc_hd__xor2_1
XFILLER_46_666 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2826 U$$3783/B1 U$$2856/A2 U$$3650/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2827/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2837 U$$2837/A U$$2839/B VGND VGND VPWR VPWR U$$2837/X sky130_fd_sc_hd__xor2_1
XFILLER_74_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2848 U$$2983/B1 U$$2866/A2 U$$2848/B1 U$$2866/B2 VGND VGND VPWR VPWR U$$2849/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_131 _290_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_21_1 U$$448/X U$$581/X U$$714/X VGND VGND VPWR VPWR dadda_fa_4_22_0/CIN
+ dadda_fa_4_21_2/A sky130_fd_sc_hd__fa_1
XFILLER_45_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2859 U$$2859/A U$$2861/B VGND VGND VPWR VPWR U$$2859/X sky130_fd_sc_hd__xor2_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_153 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 _183_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_426_ _431_/CLK _426_/D VGND VGND VPWR VPWR _426_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_197 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4407_1782 VGND VGND VPWR VPWR U$$4407_1782/HI U$$4407/B sky130_fd_sc_hd__conb_1
XFILLER_186_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_357_ _486_/CLK _357_/D VGND VGND VPWR VPWR _357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_288_ _526_/CLK _288_/D VGND VGND VPWR VPWR _288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_80_5 dadda_fa_2_80_5/A dadda_fa_2_80_5/B dadda_fa_2_80_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_2/A dadda_fa_4_80_0/A sky130_fd_sc_hd__fa_2
XFILLER_5_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_73_4 dadda_fa_2_73_4/A dadda_fa_2_73_4/B dadda_fa_2_73_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/CIN dadda_fa_3_73_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_66_3 dadda_fa_2_66_3/A dadda_fa_2_66_3/B dadda_fa_2_66_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/B dadda_fa_3_66_3/B sky130_fd_sc_hd__fa_1
XFILLER_57_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_59_2 dadda_fa_2_59_2/A dadda_fa_2_59_2/B dadda_fa_2_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/A dadda_fa_3_59_3/A sky130_fd_sc_hd__fa_1
XFILLER_110_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 a[12] VGND VGND VPWR VPWR _628_/D sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_5_36_1 dadda_fa_5_36_1/A dadda_fa_5_36_1/B dadda_fa_5_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_37_0/B dadda_fa_7_36_0/A sky130_fd_sc_hd__fa_1
XFILLER_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_29_0 dadda_fa_5_29_0/A dadda_fa_5_29_0/B dadda_fa_5_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_30_0/A dadda_fa_6_29_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_110_1 dadda_fa_5_110_1/A dadda_fa_5_110_1/B dadda_fa_5_110_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_111_0/B dadda_fa_7_110_0/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$2 _426_/Q _298_/Q VGND VGND VPWR VPWR final_adder.U$$497/B1 final_adder.U$$624/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_5_103_0 dadda_fa_5_103_0/A dadda_fa_5_103_0/B dadda_fa_5_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_104_0/A dadda_fa_6_103_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_161_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput330 _218_/Q VGND VGND VPWR VPWR o[50] sky130_fd_sc_hd__buf_2
Xoutput341 _228_/Q VGND VGND VPWR VPWR o[60] sky130_fd_sc_hd__buf_2
XFILLER_156_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput352 _238_/Q VGND VGND VPWR VPWR o[70] sky130_fd_sc_hd__buf_2
XFILLER_0_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput363 _248_/Q VGND VGND VPWR VPWR o[80] sky130_fd_sc_hd__buf_2
XFILLER_160_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput374 _258_/Q VGND VGND VPWR VPWR o[90] sky130_fd_sc_hd__buf_2
XFILLER_82_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_2 U$$2789/X U$$2922/X U$$3055/X VGND VGND VPWR VPWR dadda_fa_2_62_1/A
+ dadda_fa_2_61_4/A sky130_fd_sc_hd__fa_1
XFILLER_56_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_54_1 U$$1179/X U$$1312/X U$$1445/X VGND VGND VPWR VPWR dadda_fa_2_55_0/CIN
+ dadda_fa_2_54_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_31_0 dadda_fa_4_31_0/A dadda_fa_4_31_0/B dadda_fa_4_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/A dadda_fa_5_31_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_47_0 U$$101/X U$$234/X U$$367/X VGND VGND VPWR VPWR dadda_fa_2_48_1/B
+ dadda_fa_2_47_4/A sky130_fd_sc_hd__fa_1
XFILLER_76_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_211_ _213_/CLK _211_/D VGND VGND VPWR VPWR _211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_894 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_83_3 dadda_fa_3_83_3/A dadda_fa_3_83_3/B dadda_fa_3_83_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_1/B dadda_fa_4_83_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_76_2 dadda_fa_3_76_2/A dadda_fa_3_76_2/B dadda_fa_3_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_1/A dadda_fa_4_76_2/B sky130_fd_sc_hd__fa_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4437_1797 VGND VGND VPWR VPWR U$$4437_1797/HI U$$4437/B sky130_fd_sc_hd__conb_1
Xdadda_fa_3_69_1 dadda_fa_3_69_1/A dadda_fa_3_69_1/B dadda_fa_3_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_0/CIN dadda_fa_4_69_2/A sky130_fd_sc_hd__fa_1
XFILLER_78_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_46_0 dadda_fa_6_46_0/A dadda_fa_6_46_0/B dadda_fa_6_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_47_0/B dadda_fa_7_46_0/CIN sky130_fd_sc_hd__fa_1
XU$$4003 U$$4003/A1 U$$4035/A2 U$$4140/B1 U$$4081/B2 VGND VGND VPWR VPWR U$$4004/A
+ sky130_fd_sc_hd__a22o_1
XU$$4014 U$$4014/A U$$4058/B VGND VGND VPWR VPWR U$$4014/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4025 U$$4160/B1 U$$4065/A2 U$$4027/A1 U$$4065/B2 VGND VGND VPWR VPWR U$$4026/A
+ sky130_fd_sc_hd__a22o_1
XU$$4036 U$$4036/A U$$4036/B VGND VGND VPWR VPWR U$$4036/X sky130_fd_sc_hd__xor2_1
XU$$3302 U$$3713/A1 U$$3356/A2 U$$3578/A1 U$$3356/B2 VGND VGND VPWR VPWR U$$3303/A
+ sky130_fd_sc_hd__a22o_1
XU$$4047 U$$4456/B1 U$$4061/A2 U$$4323/A1 U$$4061/B2 VGND VGND VPWR VPWR U$$4048/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4058 U$$4058/A U$$4058/B VGND VGND VPWR VPWR U$$4058/X sky130_fd_sc_hd__xor2_1
XFILLER_93_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3313 U$$3313/A U$$3363/B VGND VGND VPWR VPWR U$$3313/X sky130_fd_sc_hd__xor2_1
XU$$3324 U$$3735/A1 U$$3368/A2 U$$3735/B1 U$$3368/B2 VGND VGND VPWR VPWR U$$3325/A
+ sky130_fd_sc_hd__a22o_1
XU$$4069 _596_/Q U$$4071/A2 U$$4206/B1 U$$4071/B2 VGND VGND VPWR VPWR U$$4070/A sky130_fd_sc_hd__a22o_1
XU$$3335 U$$3335/A U$$3369/B VGND VGND VPWR VPWR U$$3335/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3346 U$$3346/A1 U$$3356/A2 _578_/Q U$$3356/B2 VGND VGND VPWR VPWR U$$3347/A sky130_fd_sc_hd__a22o_1
XU$$2601 U$$2601/A U$$2603/A VGND VGND VPWR VPWR U$$2601/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2612 U$$2612/A U$$2698/B VGND VGND VPWR VPWR U$$2612/X sky130_fd_sc_hd__xor2_1
XFILLER_206_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3357 U$$3357/A U$$3357/B VGND VGND VPWR VPWR U$$3357/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_105_2 dadda_fa_4_105_2/A dadda_fa_4_105_2/B dadda_fa_4_105_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/CIN dadda_fa_5_105_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_185_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3368 U$$3642/A1 U$$3368/A2 U$$3505/B1 U$$3368/B2 VGND VGND VPWR VPWR U$$3369/A
+ sky130_fd_sc_hd__a22o_1
XU$$2623 U$$3717/B1 U$$2653/A2 U$$2625/A1 U$$2653/B2 VGND VGND VPWR VPWR U$$2624/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2634 U$$2634/A U$$2688/B VGND VGND VPWR VPWR U$$2634/X sky130_fd_sc_hd__xor2_1
XU$$3379 U$$3379/A U$$3407/B VGND VGND VPWR VPWR U$$3379/X sky130_fd_sc_hd__xor2_1
XU$$2645 U$$3876/B1 U$$2697/A2 U$$3741/B1 U$$2697/B2 VGND VGND VPWR VPWR U$$2646/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1900 U$$1900/A U$$1916/B VGND VGND VPWR VPWR U$$1900/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2656 U$$2656/A U$$2664/B VGND VGND VPWR VPWR U$$2656/X sky130_fd_sc_hd__xor2_1
XU$$1911 U$$3418/A1 U$$1915/A2 U$$678/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1912/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2667 U$$4035/B1 U$$2705/A2 U$$3902/A1 U$$2705/B2 VGND VGND VPWR VPWR U$$2668/A
+ sky130_fd_sc_hd__a22o_1
XU$$1922 U$$1920/Y _644_/Q _643_/Q U$$1921/X U$$1918/Y VGND VGND VPWR VPWR U$$1922/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_62_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1933 U$$1933/A U$$1983/B VGND VGND VPWR VPWR U$$1933/X sky130_fd_sc_hd__xor2_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2678 U$$2678/A U$$2708/B VGND VGND VPWR VPWR U$$2678/X sky130_fd_sc_hd__xor2_1
XU$$2689 U$$908/A1 U$$2729/A2 U$$4061/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2690/A
+ sky130_fd_sc_hd__a22o_1
XU$$1944 U$$848/A1 U$$2010/A2 U$$848/B1 U$$2010/B2 VGND VGND VPWR VPWR U$$1945/A sky130_fd_sc_hd__a22o_1
XFILLER_203_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1955 U$$1955/A U$$1957/B VGND VGND VPWR VPWR U$$1955/X sky130_fd_sc_hd__xor2_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1966 U$$2375/B1 U$$1982/A2 U$$50/A1 U$$1982/B2 VGND VGND VPWR VPWR U$$1967/A sky130_fd_sc_hd__a22o_1
XFILLER_203_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1977 U$$1977/A U$$1977/B VGND VGND VPWR VPWR U$$1977/X sky130_fd_sc_hd__xor2_1
XFILLER_15_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1988 U$$3495/A1 U$$2040/A2 U$$2947/B1 U$$2040/B2 VGND VGND VPWR VPWR U$$1989/A
+ sky130_fd_sc_hd__a22o_1
XU$$1999 U$$1999/A U$$2003/B VGND VGND VPWR VPWR U$$1999/X sky130_fd_sc_hd__xor2_1
X_409_ _538_/CLK _409_/D VGND VGND VPWR VPWR _409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_119_0 dadda_fa_7_119_0/A dadda_fa_7_119_0/B dadda_fa_7_119_0/CIN VGND
+ VGND VPWR VPWR _544_/D _415_/D sky130_fd_sc_hd__fa_1
XFILLER_179_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_947 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_71_1 dadda_fa_2_71_1/A dadda_fa_2_71_1/B dadda_fa_2_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_0/CIN dadda_fa_3_71_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_64_0 dadda_fa_2_64_0/A dadda_fa_2_64_0/B dadda_fa_2_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_0/B dadda_fa_3_64_2/B sky130_fd_sc_hd__fa_1
XFILLER_5_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater800 U$$2387/B2 VGND VGND VPWR VPWR U$$2367/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$607 ANTENNA_9/DIODE final_adder.U$$734/B final_adder.U$$607/B1 VGND
+ VGND VPWR VPWR final_adder.U$$735/B sky130_fd_sc_hd__a21o_1
Xrepeater811 U$$2274/B2 VGND VGND VPWR VPWR U$$2302/B2 sky130_fd_sc_hd__buf_6
XFILLER_97_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater822 U$$2060/X VGND VGND VPWR VPWR U$$2185/B2 sky130_fd_sc_hd__buf_6
XFILLER_56_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$629 final_adder.U$$7/SUM final_adder.U$$629/B VGND VGND VPWR VPWR
+ _175_/D sky130_fd_sc_hd__xor2_1
Xrepeater833 U$$1907/B2 VGND VGND VPWR VPWR U$$1851/B2 sky130_fd_sc_hd__buf_4
XFILLER_38_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater844 U$$1778/B2 VGND VGND VPWR VPWR U$$1768/B2 sky130_fd_sc_hd__buf_6
Xrepeater855 U$$1512/X VGND VGND VPWR VPWR U$$1607/B2 sky130_fd_sc_hd__buf_4
XFILLER_38_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater866 U$$1478/B2 VGND VGND VPWR VPWR U$$1442/B2 sky130_fd_sc_hd__buf_4
XFILLER_42_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater877 U$$1367/B2 VGND VGND VPWR VPWR U$$1355/B2 sky130_fd_sc_hd__buf_6
XFILLER_65_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater888 U$$52/B2 VGND VGND VPWR VPWR U$$8/B2 sky130_fd_sc_hd__clkbuf_4
XU$$40 U$$40/A1 U$$62/A2 U$$42/A1 U$$62/B2 VGND VGND VPWR VPWR U$$41/A sky130_fd_sc_hd__a22o_1
Xrepeater899 U$$4480/B2 VGND VGND VPWR VPWR U$$4468/B2 sky130_fd_sc_hd__buf_4
XU$$51 U$$51/A U$$99/B VGND VGND VPWR VPWR U$$51/X sky130_fd_sc_hd__xor2_1
XU$$62 U$$62/A1 U$$62/A2 U$$64/A1 U$$62/B2 VGND VGND VPWR VPWR U$$63/A sky130_fd_sc_hd__a22o_1
XU$$73 U$$73/A U$$81/B VGND VGND VPWR VPWR U$$73/X sky130_fd_sc_hd__xor2_1
XFILLER_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$84 U$$84/A1 U$$84/A2 U$$84/B1 U$$84/B2 VGND VGND VPWR VPWR U$$85/A sky130_fd_sc_hd__a22o_1
XU$$3880 U$$4154/A1 U$$3916/A2 U$$4154/B1 U$$3916/B2 VGND VGND VPWR VPWR U$$3881/A
+ sky130_fd_sc_hd__a22o_1
XU$$3891 U$$3891/A U$$3917/B VGND VGND VPWR VPWR U$$3891/X sky130_fd_sc_hd__xor2_1
XU$$95 U$$95/A U$$99/B VGND VGND VPWR VPWR U$$95/X sky130_fd_sc_hd__xor2_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_20 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _282_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_42 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_53 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_64 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_75 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_86 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_97 _287_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_4_93_2 dadda_fa_4_93_2/A dadda_fa_4_93_2/B dadda_fa_4_93_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/CIN dadda_fa_5_93_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_86_1 dadda_fa_4_86_1/A dadda_fa_4_86_1/B dadda_fa_4_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/B dadda_fa_5_86_1/B sky130_fd_sc_hd__fa_1
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_63_0 dadda_fa_7_63_0/A dadda_fa_7_63_0/B dadda_fa_7_63_0/CIN VGND VGND
+ VPWR VPWR _488_/D _359_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_79_0 dadda_fa_4_79_0/A dadda_fa_4_79_0/B dadda_fa_4_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/A dadda_fa_5_79_1/A sky130_fd_sc_hd__fa_1
XFILLER_121_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1020 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1207 U$$1207/A U$$1209/B VGND VGND VPWR VPWR U$$1207/X sky130_fd_sc_hd__xor2_1
XFILLER_46_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1218 U$$2586/B1 U$$1224/A2 U$$2588/B1 U$$1224/B2 VGND VGND VPWR VPWR U$$1219/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1229 U$$1229/A U$$1232/A VGND VGND VPWR VPWR U$$1229/X sky130_fd_sc_hd__xor2_1
XFILLER_31_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1376_1718 VGND VGND VPWR VPWR U$$1376_1718/HI U$$1376/A1 sky130_fd_sc_hd__conb_1
XFILLER_12_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_81_0 dadda_fa_3_81_0/A dadda_fa_3_81_0/B dadda_fa_3_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_0/B dadda_fa_4_81_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_194_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2335_1733 VGND VGND VPWR VPWR U$$2335_1733/HI U$$2335/A1 sky130_fd_sc_hd__conb_1
XFILLER_4_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3110 U$$3245/B1 U$$3110/A2 U$$3112/A1 U$$3110/B2 VGND VGND VPWR VPWR U$$3111/A
+ sky130_fd_sc_hd__a22o_1
XU$$3121 U$$3121/A U$$3121/B VGND VGND VPWR VPWR U$$3121/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_43_5 dadda_fa_2_43_5/A dadda_fa_2_43_5/B dadda_fa_2_43_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_2/A dadda_fa_4_43_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_4_110_0 input141/X dadda_fa_4_110_0/B dadda_fa_4_110_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_5_111_0/A dadda_fa_5_110_1/A sky130_fd_sc_hd__fa_1
XFILLER_47_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3132 U$$3132/A1 U$$3132/A2 U$$3132/B1 U$$3132/B2 VGND VGND VPWR VPWR U$$3133/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3143 U$$3143/A U$$3145/B VGND VGND VPWR VPWR U$$3143/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1060 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3154 U$$3288/A U$$3154/B VGND VGND VPWR VPWR U$$3154/X sky130_fd_sc_hd__and2_1
XU$$2420 U$$2420/A U$$2462/B VGND VGND VPWR VPWR U$$2420/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_36_4 U$$2340/X U$$2473/X U$$2517/B VGND VGND VPWR VPWR dadda_fa_3_37_1/CIN
+ dadda_fa_3_36_3/CIN sky130_fd_sc_hd__fa_1
XU$$3165 U$$3713/A1 U$$3215/A2 U$$3578/A1 U$$3215/B2 VGND VGND VPWR VPWR U$$3166/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2431 U$$785/B1 U$$2435/A2 U$$2431/B1 U$$2435/B2 VGND VGND VPWR VPWR U$$2432/A
+ sky130_fd_sc_hd__a22o_1
XU$$3176 U$$3176/A U$$3218/B VGND VGND VPWR VPWR U$$3176/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3187 U$$856/B1 U$$3209/A2 U$$3187/B1 U$$3209/B2 VGND VGND VPWR VPWR U$$3188/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2442 U$$2442/A U$$2442/B VGND VGND VPWR VPWR U$$2442/X sky130_fd_sc_hd__xor2_1
XU$$2453 _610_/Q U$$2463/A2 _611_/Q U$$2463/B2 VGND VGND VPWR VPWR U$$2454/A sky130_fd_sc_hd__a22o_1
XU$$3198 U$$3198/A U$$3236/B VGND VGND VPWR VPWR U$$3198/X sky130_fd_sc_hd__xor2_1
XU$$2464 U$$2464/A U$$2465/A VGND VGND VPWR VPWR U$$2464/X sky130_fd_sc_hd__xor2_1
XU$$2475 U$$2475/A U$$2517/B VGND VGND VPWR VPWR U$$2475/X sky130_fd_sc_hd__xor2_1
XU$$1730 U$$86/A1 U$$1736/A2 U$$88/A1 U$$1736/B2 VGND VGND VPWR VPWR U$$1731/A sky130_fd_sc_hd__a22o_1
XFILLER_34_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2486 U$$3717/B1 U$$2530/A2 U$$2625/A1 U$$2530/B2 VGND VGND VPWR VPWR U$$2487/A
+ sky130_fd_sc_hd__a22o_1
XU$$1741 U$$1741/A U$$1747/B VGND VGND VPWR VPWR U$$1741/X sky130_fd_sc_hd__xor2_1
XFILLER_72_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1752 U$$3122/A1 U$$1762/A2 U$$3124/A1 U$$1762/B2 VGND VGND VPWR VPWR U$$1753/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2497 U$$2497/A U$$2517/B VGND VGND VPWR VPWR U$$2497/X sky130_fd_sc_hd__xor2_1
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1763 U$$1763/A U$$1763/B VGND VGND VPWR VPWR U$$1763/X sky130_fd_sc_hd__xor2_1
XFILLER_210_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1774 U$$4238/B1 U$$1778/A2 U$$4105/A1 U$$1778/B2 VGND VGND VPWR VPWR U$$1775/A
+ sky130_fd_sc_hd__a22o_1
XU$$1785 U$$1783/Y _642_/Q _641_/Q U$$1784/X U$$1781/Y VGND VGND VPWR VPWR U$$1785/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_194_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1796 U$$1796/A U$$1820/B VGND VGND VPWR VPWR U$$1796/X sky130_fd_sc_hd__xor2_1
XFILLER_175_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_96_0 dadda_fa_5_96_0/A dadda_fa_5_96_0/B dadda_fa_5_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_97_0/A dadda_fa_6_96_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput40 a[45] VGND VGND VPWR VPWR _661_/D sky130_fd_sc_hd__clkbuf_1
Xinput51 a[55] VGND VGND VPWR VPWR _671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput62 a[7] VGND VGND VPWR VPWR _623_/D sky130_fd_sc_hd__clkbuf_2
Xinput73 b[17] VGND VGND VPWR VPWR _569_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput84 b[27] VGND VGND VPWR VPWR _579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput95 b[37] VGND VGND VPWR VPWR _589_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$415 final_adder.U$$332/B final_adder.U$$670/B final_adder.U$$281/X
+ VGND VGND VPWR VPWR final_adder.U$$674/B sky130_fd_sc_hd__a21o_1
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater630 U$$1345/A2 VGND VGND VPWR VPWR U$$1367/A2 sky130_fd_sc_hd__buf_6
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$437 final_adder.U$$260/B final_adder.U$$630/B final_adder.U$$137/X
+ VGND VGND VPWR VPWR final_adder.U$$632/B sky130_fd_sc_hd__a21o_1
XFILLER_84_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater641 U$$999/B2 VGND VGND VPWR VPWR U$$979/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater652 U$$924/B2 VGND VGND VPWR VPWR U$$896/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$459 final_adder.U$$282/B final_adder.U$$674/B final_adder.U$$181/X
+ VGND VGND VPWR VPWR final_adder.U$$676/B sky130_fd_sc_hd__a21o_1
Xrepeater663 U$$690/X VGND VGND VPWR VPWR U$$809/B2 sky130_fd_sc_hd__buf_6
XFILLER_84_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater674 U$$4381/B2 VGND VGND VPWR VPWR U$$4369/B2 sky130_fd_sc_hd__buf_6
XU$$309 U$$309/A U$$309/B VGND VGND VPWR VPWR U$$309/X sky130_fd_sc_hd__xor2_1
XFILLER_84_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater685 U$$545/B2 VGND VGND VPWR VPWR U$$517/B2 sky130_fd_sc_hd__buf_4
Xrepeater696 U$$4081/B2 VGND VGND VPWR VPWR U$$4105/B2 sky130_fd_sc_hd__buf_6
XFILLER_203_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_926 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1209 U$$952/A1 VGND VGND VPWR VPWR U$$950/B1 sky130_fd_sc_hd__buf_8
XU$$2874_1742 VGND VGND VPWR VPWR U$$2874_1742/HI U$$2874/B1 sky130_fd_sc_hd__conb_1
XFILLER_180_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_105_1 U$$4074/X U$$4207/X U$$4340/X VGND VGND VPWR VPWR dadda_fa_4_106_0/CIN
+ dadda_fa_4_105_2/A sky130_fd_sc_hd__fa_1
XFILLER_106_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_126_0 U$$4515/X input158/X dadda_fa_6_126_0/CIN VGND VGND VPWR VPWR dadda_fa_7_127_0/B
+ dadda_fa_7_126_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_69_4 U$$2007/X U$$2140/X U$$2273/X VGND VGND VPWR VPWR dadda_fa_1_70_7/B
+ dadda_fa_2_69_0/A sky130_fd_sc_hd__fa_1
XTAP_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_46_3 dadda_fa_3_46_3/A dadda_fa_3_46_3/B dadda_fa_3_46_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_1/B dadda_fa_4_46_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$810 U$$810/A U$$810/B VGND VGND VPWR VPWR U$$810/X sky130_fd_sc_hd__xor2_1
XU$$821 U$$821/A VGND VGND VPWR VPWR U$$821/Y sky130_fd_sc_hd__inv_1
XFILLER_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_528 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_674_ _674_/CLK _674_/D VGND VGND VPWR VPWR _674_/Q sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_3_39_2 dadda_fa_3_39_2/A dadda_fa_3_39_2/B dadda_fa_3_39_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_1/A dadda_fa_4_39_2/B sky130_fd_sc_hd__fa_1
XTAP_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$832 U$$969/A1 U$$860/A2 U$$971/A1 U$$860/B2 VGND VGND VPWR VPWR U$$833/A sky130_fd_sc_hd__a22o_1
XU$$843 U$$843/A U$$879/B VGND VGND VPWR VPWR U$$843/X sky130_fd_sc_hd__xor2_1
XFILLER_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$854 U$$854/A1 U$$924/A2 U$$993/A1 U$$924/B2 VGND VGND VPWR VPWR U$$855/A sky130_fd_sc_hd__a22o_1
XFILLER_204_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1004 U$$1004/A U$$980/B VGND VGND VPWR VPWR U$$1004/X sky130_fd_sc_hd__xor2_1
XU$$865 U$$865/A U$$925/B VGND VGND VPWR VPWR U$$865/X sky130_fd_sc_hd__xor2_1
XU$$876 U$$876/A1 U$$878/A2 U$$878/A1 U$$878/B2 VGND VGND VPWR VPWR U$$877/A sky130_fd_sc_hd__a22o_1
XFILLER_44_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1015 U$$878/A1 U$$1039/A2 U$$880/A1 U$$1039/B2 VGND VGND VPWR VPWR U$$1016/A sky130_fd_sc_hd__a22o_1
XFILLER_17_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1026 U$$1026/A U$$998/B VGND VGND VPWR VPWR U$$1026/X sky130_fd_sc_hd__xor2_1
XU$$887 U$$887/A U$$929/B VGND VGND VPWR VPWR U$$887/X sky130_fd_sc_hd__xor2_1
XFILLER_71_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1037 U$$78/A1 U$$1039/A2 U$$80/A1 U$$1039/B2 VGND VGND VPWR VPWR U$$1038/A sky130_fd_sc_hd__a22o_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$898 U$$898/A1 U$$906/A2 U$$900/A1 U$$906/B2 VGND VGND VPWR VPWR U$$899/A sky130_fd_sc_hd__a22o_1
XU$$1048 U$$1048/A U$$1090/B VGND VGND VPWR VPWR U$$1048/X sky130_fd_sc_hd__xor2_1
XFILLER_32_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1059 U$$2838/B1 U$$1065/A2 U$$2705/A1 U$$1065/B2 VGND VGND VPWR VPWR U$$1060/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_975 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_891 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1710 _552_/Q VGND VGND VPWR VPWR U$$4392/A1 sky130_fd_sc_hd__buf_6
XFILLER_171_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_675 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_41_2 U$$2350/X U$$2483/X U$$2616/X VGND VGND VPWR VPWR dadda_fa_3_42_1/A
+ dadda_fa_3_41_3/A sky130_fd_sc_hd__fa_1
XFILLER_19_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_34_1 U$$740/X U$$873/X U$$1006/X VGND VGND VPWR VPWR dadda_fa_3_35_0/CIN
+ dadda_fa_3_34_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_207_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_11_0 U$$694/X input151/X dadda_fa_5_11_0/CIN VGND VGND VPWR VPWR dadda_fa_6_12_0/A
+ dadda_fa_6_11_0/CIN sky130_fd_sc_hd__fa_1
XU$$2250 U$$467/B1 U$$2302/A2 U$$4031/B1 U$$2302/B2 VGND VGND VPWR VPWR U$$2251/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_27_0 U$$61/X U$$194/X U$$327/X VGND VGND VPWR VPWR dadda_fa_3_28_2/A dadda_fa_3_27_3/B
+ sky130_fd_sc_hd__fa_1
XU$$2261 U$$2261/A U$$2269/B VGND VGND VPWR VPWR U$$2261/X sky130_fd_sc_hd__xor2_1
XU$$2272 U$$3642/A1 U$$2274/A2 U$$3505/B1 U$$2274/B2 VGND VGND VPWR VPWR U$$2273/A
+ sky130_fd_sc_hd__a22o_1
XU$$2283 U$$2283/A U$$2299/B VGND VGND VPWR VPWR U$$2283/X sky130_fd_sc_hd__xor2_1
XU$$2294 U$$785/B1 U$$2298/A2 U$$2431/B1 U$$2298/B2 VGND VGND VPWR VPWR U$$2295/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_959 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1560 U$$1560/A U$$1598/B VGND VGND VPWR VPWR U$$1560/X sky130_fd_sc_hd__xor2_1
XU$$1571 U$$749/A1 U$$1577/A2 U$$3217/A1 U$$1577/B2 VGND VGND VPWR VPWR U$$1572/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1582 U$$1582/A U$$1628/B VGND VGND VPWR VPWR U$$1582/X sky130_fd_sc_hd__xor2_1
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1593 U$$86/A1 U$$1597/A2 U$$88/A1 U$$1597/B2 VGND VGND VPWR VPWR U$$1594/A sky130_fd_sc_hd__a22o_1
XFILLER_124_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_86_4 U$$3105/X U$$3238/X U$$3371/X VGND VGND VPWR VPWR dadda_fa_2_87_4/A
+ dadda_fa_2_86_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_79_3 U$$2293/X U$$2426/X U$$2559/X VGND VGND VPWR VPWR dadda_fa_2_80_1/B
+ dadda_fa_2_79_4/B sky130_fd_sc_hd__fa_1
XFILLER_83_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_56_2 dadda_fa_4_56_2/A dadda_fa_4_56_2/B dadda_fa_4_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/CIN dadda_fa_5_56_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_44_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$201 final_adder.U$$695/A final_adder.U$$567/B1 final_adder.U$$201/B1
+ VGND VGND VPWR VPWR final_adder.U$$201/X sky130_fd_sc_hd__a21o_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$212 final_adder.U$$707/A final_adder.U$$706/A VGND VGND VPWR VPWR
+ final_adder.U$$298/B sky130_fd_sc_hd__and2_1
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$223 final_adder.U$$717/A final_adder.U$$589/B1 final_adder.U$$223/B1
+ VGND VGND VPWR VPWR final_adder.U$$223/X sky130_fd_sc_hd__a21o_1
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_49_1 dadda_fa_4_49_1/A dadda_fa_4_49_1/B dadda_fa_4_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/B dadda_fa_5_49_1/B sky130_fd_sc_hd__fa_1
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$234 final_adder.U$$729/A final_adder.U$$728/A VGND VGND VPWR VPWR
+ final_adder.U$$308/A sky130_fd_sc_hd__and2_1
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$245 final_adder.U$$739/A final_adder.U$$611/B1 final_adder.U$$245/B1
+ VGND VGND VPWR VPWR final_adder.U$$245/X sky130_fd_sc_hd__a21o_1
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater460 U$$3968/A2 VGND VGND VPWR VPWR U$$3958/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_7_26_0 dadda_fa_7_26_0/A dadda_fa_7_26_0/B dadda_fa_7_26_0/CIN VGND VGND
+ VPWR VPWR _451_/D _322_/D sky130_fd_sc_hd__fa_1
XFILLER_45_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$106 U$$515/B1 U$$118/A2 U$$517/B1 U$$118/B2 VGND VGND VPWR VPWR U$$107/A sky130_fd_sc_hd__a22o_1
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater471 U$$3674/A2 VGND VGND VPWR VPWR U$$3628/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$267 final_adder.U$$266/A final_adder.U$$149/X final_adder.U$$151/X
+ VGND VGND VPWR VPWR final_adder.U$$267/X sky130_fd_sc_hd__a21o_1
XU$$117 U$$117/A U$$117/B VGND VGND VPWR VPWR U$$117/X sky130_fd_sc_hd__xor2_1
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater482 U$$3429/X VGND VGND VPWR VPWR U$$3537/A2 sky130_fd_sc_hd__buf_6
XFILLER_85_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$278 final_adder.U$$278/A final_adder.U$$278/B VGND VGND VPWR VPWR
+ final_adder.U$$330/A sky130_fd_sc_hd__and2_2
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$128 U$$676/A1 U$$128/A2 U$$676/B1 U$$128/B2 VGND VGND VPWR VPWR U$$129/A sky130_fd_sc_hd__a22o_1
Xrepeater493 U$$3292/X VGND VGND VPWR VPWR U$$3408/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$289 final_adder.U$$288/A final_adder.U$$193/X final_adder.U$$195/X
+ VGND VGND VPWR VPWR final_adder.U$$289/X sky130_fd_sc_hd__a21o_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$139 U$$272/B VGND VGND VPWR VPWR U$$139/Y sky130_fd_sc_hd__inv_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_390_ _520_/CLK _390_/D VGND VGND VPWR VPWR _390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_222 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1006 U$$2843/B VGND VGND VPWR VPWR U$$2839/B sky130_fd_sc_hd__buf_6
XFILLER_181_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1017 U$$2734/B VGND VGND VPWR VPWR U$$2730/B sky130_fd_sc_hd__buf_6
XFILLER_107_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1028 _653_/Q VGND VGND VPWR VPWR U$$2603/A sky130_fd_sc_hd__buf_12
Xrepeater1039 U$$2243/B VGND VGND VPWR VPWR U$$2241/B sky130_fd_sc_hd__buf_8
XFILLER_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1040 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_51_1 dadda_fa_3_51_1/A dadda_fa_3_51_1/B dadda_fa_3_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_0/CIN dadda_fa_4_51_2/A sky130_fd_sc_hd__fa_1
Xinput230 c[76] VGND VGND VPWR VPWR input230/X sky130_fd_sc_hd__clkbuf_4
Xinput241 c[86] VGND VGND VPWR VPWR input241/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_0_67_1 U$$540/X U$$673/X U$$806/X VGND VGND VPWR VPWR dadda_fa_1_68_5/CIN
+ dadda_fa_1_67_7/CIN sky130_fd_sc_hd__fa_1
Xinput252 c[96] VGND VGND VPWR VPWR input252/X sky130_fd_sc_hd__buf_4
XTAP_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_44_0 dadda_fa_3_44_0/A dadda_fa_3_44_0/B dadda_fa_3_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_0/B dadda_fa_4_44_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$640 U$$912/B1 U$$650/A2 U$$914/B1 U$$650/B2 VGND VGND VPWR VPWR U$$641/A sky130_fd_sc_hd__a22o_1
XFILLER_205_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_657_ _662_/CLK _657_/D VGND VGND VPWR VPWR _657_/Q sky130_fd_sc_hd__dfxtp_4
XU$$651 U$$651/A U$$651/B VGND VGND VPWR VPWR U$$651/X sky130_fd_sc_hd__xor2_1
XU$$662 U$$936/A1 U$$668/A2 U$$938/A1 U$$670/B2 VGND VGND VPWR VPWR U$$663/A sky130_fd_sc_hd__a22o_1
XU$$673 U$$673/A U$$685/A VGND VGND VPWR VPWR U$$673/X sky130_fd_sc_hd__xor2_1
XFILLER_44_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$684 U$$684/A VGND VGND VPWR VPWR U$$684/Y sky130_fd_sc_hd__inv_1
XU$$695 U$$695/A1 U$$725/A2 U$$695/B1 U$$725/B2 VGND VGND VPWR VPWR U$$696/A sky130_fd_sc_hd__a22o_1
X_588_ _588_/CLK _588_/D VGND VGND VPWR VPWR _588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1039 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_101_0 dadda_fa_7_101_0/A dadda_fa_7_101_0/B dadda_fa_7_101_0/CIN VGND
+ VGND VPWR VPWR _526_/D _397_/D sky130_fd_sc_hd__fa_1
XFILLER_157_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_636 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_96_3 U$$3657/X U$$3790/X U$$3923/X VGND VGND VPWR VPWR dadda_fa_3_97_1/B
+ dadda_fa_3_96_3/B sky130_fd_sc_hd__fa_1
XFILLER_144_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1540 U$$2375/B1 VGND VGND VPWR VPWR U$$48/A1 sky130_fd_sc_hd__buf_6
Xrepeater1551 U$$866/B1 VGND VGND VPWR VPWR U$$46/A1 sky130_fd_sc_hd__buf_8
Xrepeater1562 U$$4154/A1 VGND VGND VPWR VPWR U$$2508/B1 sky130_fd_sc_hd__buf_4
XFILLER_153_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_89_2 U$$4175/X U$$4308/X U$$4441/X VGND VGND VPWR VPWR dadda_fa_3_90_1/A
+ dadda_fa_3_89_3/A sky130_fd_sc_hd__fa_1
Xrepeater1573 U$$999/A1 VGND VGND VPWR VPWR U$$3054/A1 sky130_fd_sc_hd__buf_6
XFILLER_98_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1584 _567_/Q VGND VGND VPWR VPWR U$$3735/B1 sky130_fd_sc_hd__buf_6
XFILLER_63_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1595 U$$3046/B1 VGND VGND VPWR VPWR U$$582/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_66_1 dadda_fa_5_66_1/A dadda_fa_5_66_1/B dadda_fa_5_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_67_0/B dadda_fa_7_66_0/A sky130_fd_sc_hd__fa_1
XFILLER_125_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_59_0 dadda_fa_5_59_0/A dadda_fa_5_59_0/B dadda_fa_5_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_60_0/A dadda_fa_6_59_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_58_8 dadda_fa_1_58_8/A dadda_fa_1_58_8/B dadda_fa_1_58_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_59_3/A dadda_fa_3_58_0/A sky130_fd_sc_hd__fa_2
XFILLER_104_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_105_0 U$$2876/Y U$$3010/X U$$3143/X VGND VGND VPWR VPWR dadda_fa_3_106_3/A
+ dadda_fa_3_105_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2080 U$$2080/A U$$2110/B VGND VGND VPWR VPWR U$$2080/X sky130_fd_sc_hd__xor2_1
XFILLER_74_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2091 U$$856/B1 U$$2135/A2 U$$3187/B1 U$$2135/B2 VGND VGND VPWR VPWR U$$2092/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1390 U$$840/B1 U$$1458/A2 U$$568/B1 U$$1458/B2 VGND VGND VPWR VPWR U$$1391/A sky130_fd_sc_hd__a22o_1
XFILLER_195_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_439 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_91_2 U$$2716/X U$$2849/X U$$2982/X VGND VGND VPWR VPWR dadda_fa_2_92_5/A
+ dadda_fa_3_91_0/A sky130_fd_sc_hd__fa_1
XFILLER_172_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_84_1 U$$1771/X U$$1904/X U$$2037/X VGND VGND VPWR VPWR dadda_fa_2_85_2/B
+ dadda_fa_2_84_4/B sky130_fd_sc_hd__fa_1
XFILLER_104_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_61_0 dadda_fa_4_61_0/A dadda_fa_4_61_0/B dadda_fa_4_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/A dadda_fa_5_61_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_77_0 U$$1358/X U$$1491/X U$$1624/X VGND VGND VPWR VPWR dadda_fa_2_78_0/B
+ dadda_fa_2_77_3/B sky130_fd_sc_hd__fa_1
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_2_104_2 U$$3540/X U$$3673/X VGND VGND VPWR VPWR dadda_fa_3_105_3/B dadda_fa_4_104_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3709 U$$3709/A1 U$$3743/A2 _554_/Q U$$3743/B2 VGND VGND VPWR VPWR U$$3710/A sky130_fd_sc_hd__a22o_1
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_675 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_302 _235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_511_ _560_/CLK _511_/D VGND VGND VPWR VPWR _511_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_313 _237_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 _238_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_335 _177_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 U$$3096/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ _442_/CLK _442_/D VGND VGND VPWR VPWR _442_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_357 _619_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_368 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_379 U$$4357/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_373_ _503_/CLK _373_/D VGND VGND VPWR VPWR _373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_99_1 dadda_fa_3_99_1/A dadda_fa_3_99_1/B dadda_fa_3_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_0/CIN dadda_fa_4_99_2/A sky130_fd_sc_hd__fa_1
XU$$3568_1753 VGND VGND VPWR VPWR U$$3568_1753/HI U$$3568/A1 sky130_fd_sc_hd__conb_1
XFILLER_142_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_76_0 dadda_fa_6_76_0/A dadda_fa_6_76_0/B dadda_fa_6_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_77_0/B dadda_fa_7_76_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_142_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_306 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$470 U$$470/A U$$484/B VGND VGND VPWR VPWR U$$470/X sky130_fd_sc_hd__xor2_1
XFILLER_63_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$481 U$$70/A1 U$$483/A2 U$$72/A1 U$$483/B2 VGND VGND VPWR VPWR U$$482/A sky130_fd_sc_hd__a22o_1
XFILLER_205_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$492 U$$492/A U$$536/B VGND VGND VPWR VPWR U$$492/X sky130_fd_sc_hd__xor2_1
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_580 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_94_0 U$$2722/X U$$2855/X U$$2988/X VGND VGND VPWR VPWR dadda_fa_3_95_0/B
+ dadda_fa_3_94_2/B sky130_fd_sc_hd__fa_1
XFILLER_145_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1370 _594_/Q VGND VGND VPWR VPWR U$$4337/B1 sky130_fd_sc_hd__buf_6
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1381 U$$2963/B1 VGND VGND VPWR VPWR U$$88/A1 sky130_fd_sc_hd__buf_4
XFILLER_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1392 U$$4470/A1 VGND VGND VPWR VPWR U$$3374/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_119_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_70_7 dadda_fa_1_70_7/A dadda_fa_1_70_7/B dadda_fa_1_70_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_2/CIN dadda_fa_2_70_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_63_6 dadda_fa_1_63_6/A dadda_fa_1_63_6/B dadda_fa_1_63_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_2/B dadda_fa_2_63_5/B sky130_fd_sc_hd__fa_1
XFILLER_68_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_56_5 U$$3178/X U$$3311/X U$$3444/X VGND VGND VPWR VPWR dadda_fa_2_57_2/A
+ dadda_fa_2_56_5/A sky130_fd_sc_hd__fa_1
XFILLER_39_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4465_1811 VGND VGND VPWR VPWR U$$4465_1811/HI U$$4465/B sky130_fd_sc_hd__conb_1
XFILLER_131_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_49_4 U$$1701/X U$$1834/X U$$1967/X VGND VGND VPWR VPWR dadda_fa_2_50_2/A
+ dadda_fa_2_49_5/A sky130_fd_sc_hd__fa_1
XFILLER_55_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_2 dadda_fa_4_19_2/A dadda_fa_4_19_2/B dadda_ha_3_19_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_20_0/CIN dadda_fa_5_19_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_93_0 dadda_fa_7_93_0/A dadda_fa_7_93_0/B dadda_fa_7_93_0/CIN VGND VGND
+ VPWR VPWR _518_/D _389_/D sky130_fd_sc_hd__fa_2
XFILLER_206_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2472_1735 VGND VGND VPWR VPWR U$$2472_1735/HI U$$2472/A1 sky130_fd_sc_hd__conb_1
XFILLER_172_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4207 U$$4207/A U$$4247/A VGND VGND VPWR VPWR U$$4207/X sky130_fd_sc_hd__xor2_1
XU$$4218 U$$4218/A1 U$$4244/A2 U$$4355/B1 U$$4244/B2 VGND VGND VPWR VPWR U$$4219/A
+ sky130_fd_sc_hd__a22o_1
XU$$4229 U$$4229/A U$$4239/B VGND VGND VPWR VPWR U$$4229/X sky130_fd_sc_hd__xor2_1
XFILLER_58_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3506 U$$3506/A U$$3506/B VGND VGND VPWR VPWR U$$3506/X sky130_fd_sc_hd__xor2_1
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3517 U$$3789/B1 U$$3519/A2 U$$3791/B1 U$$3519/B2 VGND VGND VPWR VPWR U$$3518/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3528 U$$3528/A U$$3538/B VGND VGND VPWR VPWR U$$3528/X sky130_fd_sc_hd__xor2_1
XFILLER_65_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3539 U$$3539/A1 U$$3429/X U$$4087/B1 U$$3430/X VGND VGND VPWR VPWR U$$3540/A sky130_fd_sc_hd__a22o_1
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2805 U$$2805/A U$$2839/B VGND VGND VPWR VPWR U$$2805/X sky130_fd_sc_hd__xor2_1
XFILLER_85_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_426 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2816 U$$4186/A1 U$$2856/A2 U$$4051/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2817/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2827 U$$2827/A U$$2827/B VGND VGND VPWR VPWR U$$2827/X sky130_fd_sc_hd__xor2_1
XFILLER_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 _179_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2838 U$$2838/A1 U$$2744/X U$$2838/B1 U$$2745/X VGND VGND VPWR VPWR U$$2839/A sky130_fd_sc_hd__a22o_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 _290_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2849 U$$2849/A U$$2875/B VGND VGND VPWR VPWR U$$2849/X sky130_fd_sc_hd__xor2_1
XANTENNA_143 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_3_21_2 U$$847/X U$$980/X U$$1113/X VGND VGND VPWR VPWR dadda_fa_4_22_1/A
+ dadda_fa_4_21_2/B sky130_fd_sc_hd__fa_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _183_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_176 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_187 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_425_ _431_/CLK _425_/D VGND VGND VPWR VPWR _425_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_198 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_356_ _485_/CLK _356_/D VGND VGND VPWR VPWR _356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_287_ _526_/CLK _287_/D VGND VGND VPWR VPWR _287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_399 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_411 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_73_5 dadda_fa_2_73_5/A dadda_fa_2_73_5/B dadda_fa_2_73_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_2/A dadda_fa_4_73_0/A sky130_fd_sc_hd__fa_1
XFILLER_151_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_66_4 dadda_fa_2_66_4/A dadda_fa_2_66_4/B dadda_fa_2_66_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/CIN dadda_fa_3_66_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_59_3 dadda_fa_2_59_3/A dadda_fa_2_59_3/B dadda_fa_2_59_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/B dadda_fa_3_59_3/B sky130_fd_sc_hd__fa_1
XFILLER_96_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 a[13] VGND VGND VPWR VPWR _629_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_5_29_1 dadda_fa_5_29_1/A dadda_fa_5_29_1/B dadda_fa_5_29_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_30_0/B dadda_fa_7_29_0/A sky130_fd_sc_hd__fa_2
XFILLER_209_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_250 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4495_1826 VGND VGND VPWR VPWR U$$4495_1826/HI U$$4495/B sky130_fd_sc_hd__conb_1
XFILLER_177_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$3 _427_/Q _299_/Q VGND VGND VPWR VPWR final_adder.U$$3/COUT final_adder.U$$625/A
+ sky130_fd_sc_hd__ha_1
XFILLER_195_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_103_1 dadda_fa_5_103_1/A dadda_fa_5_103_1/B dadda_fa_5_103_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_104_0/B dadda_fa_7_103_0/A sky130_fd_sc_hd__fa_1
XFILLER_118_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput320 _209_/Q VGND VGND VPWR VPWR o[41] sky130_fd_sc_hd__buf_2
Xoutput331 _219_/Q VGND VGND VPWR VPWR o[51] sky130_fd_sc_hd__buf_2
XFILLER_160_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput342 _229_/Q VGND VGND VPWR VPWR o[61] sky130_fd_sc_hd__buf_2
Xoutput353 _239_/Q VGND VGND VPWR VPWR o[71] sky130_fd_sc_hd__buf_2
XFILLER_156_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput364 _249_/Q VGND VGND VPWR VPWR o[81] sky130_fd_sc_hd__buf_2
XFILLER_126_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput375 _259_/Q VGND VGND VPWR VPWR o[91] sky130_fd_sc_hd__buf_2
XFILLER_142_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_3 U$$3188/X U$$3321/X U$$3454/X VGND VGND VPWR VPWR dadda_fa_2_62_1/B
+ dadda_fa_2_61_4/B sky130_fd_sc_hd__fa_1
XFILLER_87_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_2 U$$1578/X U$$1711/X U$$1844/X VGND VGND VPWR VPWR dadda_fa_2_55_1/A
+ dadda_fa_2_54_4/A sky130_fd_sc_hd__fa_1
XFILLER_142_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_31_1 dadda_fa_4_31_1/A dadda_fa_4_31_1/B dadda_fa_4_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/B dadda_fa_5_31_1/B sky130_fd_sc_hd__fa_1
XFILLER_132_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_47_1 U$$500/X U$$633/X U$$766/X VGND VGND VPWR VPWR dadda_fa_2_48_1/CIN
+ dadda_fa_2_47_4/B sky130_fd_sc_hd__fa_1
XFILLER_71_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_24_0 dadda_fa_4_24_0/A dadda_fa_4_24_0/B dadda_fa_4_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/A dadda_fa_5_24_1/A sky130_fd_sc_hd__fa_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_210_ _213_/CLK _210_/D VGND VGND VPWR VPWR _210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_926 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_76_3 dadda_fa_3_76_3/A dadda_fa_3_76_3/B dadda_fa_3_76_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_1/B dadda_fa_4_76_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_69_2 dadda_fa_3_69_2/A dadda_fa_3_69_2/B dadda_fa_3_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_1/A dadda_fa_4_69_2/B sky130_fd_sc_hd__fa_1
XFILLER_78_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4004 U$$4004/A U$$4036/B VGND VGND VPWR VPWR U$$4004/X sky130_fd_sc_hd__xor2_1
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4015 _569_/Q U$$4029/A2 U$$4154/A1 U$$4029/B2 VGND VGND VPWR VPWR U$$4016/A sky130_fd_sc_hd__a22o_1
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4026 U$$4026/A U$$4044/B VGND VGND VPWR VPWR U$$4026/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_39_0 dadda_fa_6_39_0/A dadda_fa_6_39_0/B dadda_fa_6_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_40_0/B dadda_fa_7_39_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4037 U$$4446/B1 U$$4095/A2 U$$4176/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4038/A
+ sky130_fd_sc_hd__a22o_1
XU$$3303 U$$3303/A U$$3357/B VGND VGND VPWR VPWR U$$3303/X sky130_fd_sc_hd__xor2_1
XU$$4048 U$$4048/A U$$4070/B VGND VGND VPWR VPWR U$$4048/X sky130_fd_sc_hd__xor2_1
XU$$4059 _591_/Q U$$4061/A2 U$$4333/B1 U$$4061/B2 VGND VGND VPWR VPWR U$$4060/A sky130_fd_sc_hd__a22o_1
XU$$3314 U$$3451/A1 U$$3320/A2 U$$3453/A1 U$$3320/B2 VGND VGND VPWR VPWR U$$3315/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3325 U$$3325/A U$$3369/B VGND VGND VPWR VPWR U$$3325/X sky130_fd_sc_hd__xor2_1
XU$$3336 U$$4432/A1 U$$3418/A2 U$$4434/A1 U$$3418/B2 VGND VGND VPWR VPWR U$$3337/A
+ sky130_fd_sc_hd__a22o_1
XU$$3347 U$$3347/A U$$3357/B VGND VGND VPWR VPWR U$$3347/X sky130_fd_sc_hd__xor2_1
XU$$2602 U$$2603/A VGND VGND VPWR VPWR U$$2602/Y sky130_fd_sc_hd__inv_1
XU$$3358 U$$3358/A1 U$$3378/A2 U$$4317/B1 U$$3378/B2 VGND VGND VPWR VPWR U$$3359/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2613 U$$556/B1 U$$2653/A2 U$$2613/B1 U$$2653/B2 VGND VGND VPWR VPWR U$$2614/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3369 U$$3369/A U$$3369/B VGND VGND VPWR VPWR U$$3369/X sky130_fd_sc_hd__xor2_1
XFILLER_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2624 U$$2624/A U$$2654/B VGND VGND VPWR VPWR U$$2624/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2635 U$$2909/A1 U$$2687/A2 U$$2909/B1 U$$2687/B2 VGND VGND VPWR VPWR U$$2636/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1901 U$$3132/B1 U$$1909/A2 U$$944/A1 U$$1909/B2 VGND VGND VPWR VPWR U$$1902/A
+ sky130_fd_sc_hd__a22o_1
XU$$2646 U$$2646/A U$$2698/B VGND VGND VPWR VPWR U$$2646/X sky130_fd_sc_hd__xor2_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2657 U$$463/B1 U$$2663/A2 U$$330/A1 U$$2663/B2 VGND VGND VPWR VPWR U$$2658/A sky130_fd_sc_hd__a22o_1
XU$$1912 U$$1912/A U$$1916/B VGND VGND VPWR VPWR U$$1912/X sky130_fd_sc_hd__xor2_1
XU$$2668 U$$2668/A U$$2706/B VGND VGND VPWR VPWR U$$2668/X sky130_fd_sc_hd__xor2_1
XU$$1923 U$$1921/B _643_/Q _644_/Q U$$1918/Y VGND VGND VPWR VPWR U$$1923/X sky130_fd_sc_hd__a22o_4
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1934 U$$2345/A1 U$$1976/A2 U$$2895/A1 U$$1976/B2 VGND VGND VPWR VPWR U$$1935/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2679 U$$3362/B1 U$$2697/A2 U$$3229/A1 U$$2697/B2 VGND VGND VPWR VPWR U$$2680/A
+ sky130_fd_sc_hd__a22o_1
XU$$1945 U$$1945/A U$$2011/B VGND VGND VPWR VPWR U$$1945/X sky130_fd_sc_hd__xor2_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1956 U$$997/A1 U$$1956/A2 U$$999/A1 U$$1956/B2 VGND VGND VPWR VPWR U$$1957/A sky130_fd_sc_hd__a22o_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1967 U$$1967/A U$$1983/B VGND VGND VPWR VPWR U$$1967/X sky130_fd_sc_hd__xor2_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1978 U$$3485/A1 U$$2028/A2 U$$3624/A1 U$$2028/B2 VGND VGND VPWR VPWR U$$1979/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_974 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_408_ _538_/CLK _408_/D VGND VGND VPWR VPWR _408_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1989 U$$1989/A U$$2043/B VGND VGND VPWR VPWR U$$1989/X sky130_fd_sc_hd__xor2_1
XFILLER_109_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_339_ _466_/CLK _339_/D VGND VGND VPWR VPWR _339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_71_2 dadda_fa_2_71_2/A dadda_fa_2_71_2/B dadda_fa_2_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/A dadda_fa_3_71_3/A sky130_fd_sc_hd__fa_2
XFILLER_29_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_100_0_1862 VGND VGND VPWR VPWR dadda_fa_2_100_0/A dadda_fa_2_100_0_1862/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_69_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_64_1 dadda_fa_2_64_1/A dadda_fa_2_64_1/B dadda_fa_2_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_0/CIN dadda_fa_3_64_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_111_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater801 U$$2395/B2 VGND VGND VPWR VPWR U$$2387/B2 sky130_fd_sc_hd__buf_6
XFILLER_29_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater812 U$$2197/X VGND VGND VPWR VPWR U$$2274/B2 sky130_fd_sc_hd__buf_4
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$619 final_adder.U$$746/A final_adder.U$$746/B final_adder.U$$619/B1
+ VGND VGND VPWR VPWR final_adder.U$$747/B sky130_fd_sc_hd__a21o_1
Xrepeater823 U$$2040/B2 VGND VGND VPWR VPWR U$$1956/B2 sky130_fd_sc_hd__buf_6
XFILLER_57_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_41_0 dadda_fa_5_41_0/A dadda_fa_5_41_0/B dadda_fa_5_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_42_0/A dadda_fa_6_41_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_57_0 dadda_fa_2_57_0/A dadda_fa_2_57_0/B dadda_fa_2_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_0/B dadda_fa_3_57_2/B sky130_fd_sc_hd__fa_1
Xrepeater834 U$$1907/B2 VGND VGND VPWR VPWR U$$1855/B2 sky130_fd_sc_hd__buf_8
Xrepeater845 U$$1778/B2 VGND VGND VPWR VPWR U$$1740/B2 sky130_fd_sc_hd__buf_12
Xrepeater856 U$$219/B2 VGND VGND VPWR VPWR U$$175/B2 sky130_fd_sc_hd__buf_6
Xrepeater867 U$$1478/B2 VGND VGND VPWR VPWR U$$1428/B2 sky130_fd_sc_hd__buf_6
Xrepeater878 U$$1345/B2 VGND VGND VPWR VPWR U$$1367/B2 sky130_fd_sc_hd__buf_6
XU$$30 U$$30/A1 U$$68/A2 U$$32/A1 U$$68/B2 VGND VGND VPWR VPWR U$$31/A sky130_fd_sc_hd__a22o_1
Xrepeater889 U$$68/B2 VGND VGND VPWR VPWR U$$52/B2 sky130_fd_sc_hd__buf_4
XU$$41 U$$41/A U$$3/A VGND VGND VPWR VPWR U$$41/X sky130_fd_sc_hd__xor2_1
XFILLER_65_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$52 U$$52/A1 U$$52/A2 U$$52/B1 U$$52/B2 VGND VGND VPWR VPWR U$$53/A sky130_fd_sc_hd__a22o_1
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$63 U$$63/A U$$3/A VGND VGND VPWR VPWR U$$63/X sky130_fd_sc_hd__xor2_1
XFILLER_37_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$74 U$$74/A1 U$$84/A2 U$$76/A1 U$$84/B2 VGND VGND VPWR VPWR U$$75/A sky130_fd_sc_hd__a22o_1
XU$$3870 U$$4007/A1 U$$3874/A2 _566_/Q U$$3874/B2 VGND VGND VPWR VPWR U$$3871/A sky130_fd_sc_hd__a22o_1
XU$$85 U$$85/A U$$85/B VGND VGND VPWR VPWR U$$85/X sky130_fd_sc_hd__xor2_1
XU$$3881 U$$3881/A U$$3917/B VGND VGND VPWR VPWR U$$3881/X sky130_fd_sc_hd__xor2_1
XU$$96 U$$96/A1 U$$98/A2 U$$98/A1 U$$98/B2 VGND VGND VPWR VPWR U$$97/A sky130_fd_sc_hd__a22o_1
XU$$3892 U$$4440/A1 U$$3910/A2 U$$4442/A1 U$$3910/B2 VGND VGND VPWR VPWR U$$3893/A
+ sky130_fd_sc_hd__a22o_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_10 ANTENNA_10/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_21 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _282_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_54 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_65 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_386 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_76 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_98 _287_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_88_0_1858 VGND VGND VPWR VPWR dadda_fa_1_88_0/A dadda_fa_1_88_0_1858/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_192_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_86_2 dadda_fa_4_86_2/A dadda_fa_4_86_2/B dadda_fa_4_86_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/CIN dadda_fa_5_86_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_79_1 dadda_fa_4_79_1/A dadda_fa_4_79_1/B dadda_fa_4_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/B dadda_fa_5_79_1/B sky130_fd_sc_hd__fa_1
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_56_0 dadda_fa_7_56_0/A dadda_fa_7_56_0/B dadda_fa_7_56_0/CIN VGND VGND
+ VPWR VPWR _481_/D _352_/D sky130_fd_sc_hd__fa_1
XFILLER_161_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1208 U$$658/B1 U$$1208/A2 U$$4224/A1 U$$1208/B2 VGND VGND VPWR VPWR U$$1209/A
+ sky130_fd_sc_hd__a22o_1
XU$$1219 U$$1219/A U$$1225/B VGND VGND VPWR VPWR U$$1219/X sky130_fd_sc_hd__xor2_1
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_667 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_81_1 dadda_fa_3_81_1/A dadda_fa_3_81_1/B dadda_fa_3_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_0/CIN dadda_fa_4_81_2/A sky130_fd_sc_hd__fa_1
XFILLER_124_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_74_0 dadda_fa_3_74_0/A dadda_fa_3_74_0/B dadda_fa_3_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_0/B dadda_fa_4_74_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_152_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3100 U$$3374/A1 U$$3144/A2 U$$4472/A1 U$$3144/B2 VGND VGND VPWR VPWR U$$3101/A
+ sky130_fd_sc_hd__a22o_1
XU$$3111 U$$3111/A U$$3111/B VGND VGND VPWR VPWR U$$3111/X sky130_fd_sc_hd__xor2_1
XU$$3122 U$$3122/A1 U$$3132/A2 U$$3124/A1 U$$3132/B2 VGND VGND VPWR VPWR U$$3123/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_110_1 dadda_fa_4_110_1/A dadda_fa_4_110_1/B dadda_fa_4_110_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_111_0/B dadda_fa_5_110_1/B sky130_fd_sc_hd__fa_1
XU$$3133 U$$3133/A U$$3133/B VGND VGND VPWR VPWR U$$3133/X sky130_fd_sc_hd__xor2_1
XFILLER_53_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3144 U$$3281/A1 U$$3144/A2 U$$3283/A1 U$$3144/B2 VGND VGND VPWR VPWR U$$3145/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_36_5 input186/X dadda_fa_2_36_5/B dadda_fa_2_36_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_37_2/A dadda_fa_4_36_0/A sky130_fd_sc_hd__fa_2
XU$$3155 U$$3153/Y _662_/Q _661_/Q U$$3154/X U$$3151/Y VGND VGND VPWR VPWR U$$3155/X
+ sky130_fd_sc_hd__a32o_1
XU$$2410 U$$2410/A U$$2436/B VGND VGND VPWR VPWR U$$2410/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1072 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2421 U$$914/A1 U$$2423/A2 U$$916/A1 U$$2423/B2 VGND VGND VPWR VPWR U$$2422/A sky130_fd_sc_hd__a22o_1
XU$$3166 U$$3166/A U$$3218/B VGND VGND VPWR VPWR U$$3166/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_103_0 dadda_fa_4_103_0/A dadda_fa_4_103_0/B dadda_fa_4_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/A dadda_fa_5_103_1/A sky130_fd_sc_hd__fa_1
XU$$3177 U$$3312/B1 U$$3231/A2 U$$4273/B1 U$$3231/B2 VGND VGND VPWR VPWR U$$3178/A
+ sky130_fd_sc_hd__a22o_1
XU$$2432 U$$2432/A U$$2436/B VGND VGND VPWR VPWR U$$2432/X sky130_fd_sc_hd__xor2_1
XU$$3188 U$$3188/A U$$3208/B VGND VGND VPWR VPWR U$$3188/X sky130_fd_sc_hd__xor2_1
XU$$2443 U$$4087/A1 U$$2451/A2 U$$4087/B1 U$$2451/B2 VGND VGND VPWR VPWR U$$2444/A
+ sky130_fd_sc_hd__a22o_1
XU$$2454 U$$2454/A U$$2465/A VGND VGND VPWR VPWR U$$2454/X sky130_fd_sc_hd__xor2_1
XU$$3199 U$$4432/A1 U$$3235/A2 U$$4434/A1 U$$3235/B2 VGND VGND VPWR VPWR U$$3200/A
+ sky130_fd_sc_hd__a22o_1
XU$$1720 U$$896/B1 U$$1768/A2 U$$761/B1 U$$1768/B2 VGND VGND VPWR VPWR U$$1721/A sky130_fd_sc_hd__a22o_1
XU$$2465 U$$2465/A VGND VGND VPWR VPWR U$$2465/Y sky130_fd_sc_hd__inv_1
XFILLER_61_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1731 U$$1731/A U$$1737/B VGND VGND VPWR VPWR U$$1731/X sky130_fd_sc_hd__xor2_1
XFILLER_61_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2476 U$$2611/B1 U$$2516/A2 U$$2478/A1 U$$2516/B2 VGND VGND VPWR VPWR U$$2477/A
+ sky130_fd_sc_hd__a22o_1
XU$$2487 U$$2487/A U$$2531/B VGND VGND VPWR VPWR U$$2487/X sky130_fd_sc_hd__xor2_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1742 U$$3112/A1 U$$1778/A2 U$$922/A1 U$$1778/B2 VGND VGND VPWR VPWR U$$1743/A
+ sky130_fd_sc_hd__a22o_1
XU$$1753 U$$1753/A U$$1763/B VGND VGND VPWR VPWR U$$1753/X sky130_fd_sc_hd__xor2_1
XU$$2498 U$$3181/B1 U$$2516/A2 U$$3046/B1 U$$2516/B2 VGND VGND VPWR VPWR U$$2499/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1764 U$$3132/B1 U$$1768/A2 U$$2586/B1 U$$1768/B2 VGND VGND VPWR VPWR U$$1765/A
+ sky130_fd_sc_hd__a22o_1
XU$$1775 U$$1775/A U$$1780/A VGND VGND VPWR VPWR U$$1775/X sky130_fd_sc_hd__xor2_1
XFILLER_43_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1786 U$$1784/B _641_/Q _642_/Q U$$1781/Y VGND VGND VPWR VPWR U$$1786/X sky130_fd_sc_hd__a22o_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1797 U$$2756/A1 U$$1859/A2 U$$2756/B1 U$$1859/B2 VGND VGND VPWR VPWR U$$1798/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_96_1 dadda_fa_5_96_1/A dadda_fa_5_96_1/B dadda_fa_5_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_97_0/B dadda_fa_7_96_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_0_76_0_1853 VGND VGND VPWR VPWR dadda_fa_0_76_0/A dadda_fa_0_76_0_1853/LO
+ sky130_fd_sc_hd__conb_1
Xinput30 a[36] VGND VGND VPWR VPWR _652_/D sky130_fd_sc_hd__clkbuf_1
Xinput41 a[46] VGND VGND VPWR VPWR _662_/D sky130_fd_sc_hd__clkbuf_1
Xinput52 a[56] VGND VGND VPWR VPWR _672_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput63 a[8] VGND VGND VPWR VPWR _624_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_200_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_89_0 dadda_fa_5_89_0/A dadda_fa_5_89_0/B dadda_fa_5_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_90_0/A dadda_fa_6_89_0/CIN sky130_fd_sc_hd__fa_1
Xinput74 b[18] VGND VGND VPWR VPWR _570_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 b[28] VGND VGND VPWR VPWR _580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput96 b[38] VGND VGND VPWR VPWR _590_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_951 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$405 final_adder.U$$322/B final_adder.U$$630/B final_adder.U$$261/X
+ VGND VGND VPWR VPWR final_adder.U$$634/B sky130_fd_sc_hd__a21o_2
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater620 U$$1500/A2 VGND VGND VPWR VPWR U$$1486/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$427 final_adder.U$$344/B final_adder.U$$718/B final_adder.U$$305/X
+ VGND VGND VPWR VPWR final_adder.U$$722/B sky130_fd_sc_hd__a21o_1
Xrepeater631 U$$1237/X VGND VGND VPWR VPWR U$$1345/A2 sky130_fd_sc_hd__buf_6
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater642 U$$999/B2 VGND VGND VPWR VPWR U$$1039/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$449 final_adder.U$$272/B final_adder.U$$654/B final_adder.U$$161/X
+ VGND VGND VPWR VPWR final_adder.U$$656/B sky130_fd_sc_hd__a21o_1
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater653 U$$948/B2 VGND VGND VPWR VPWR U$$924/B2 sky130_fd_sc_hd__buf_6
Xrepeater664 U$$622/B2 VGND VGND VPWR VPWR U$$574/B2 sky130_fd_sc_hd__buf_4
XFILLER_42_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater675 U$$4345/B2 VGND VGND VPWR VPWR U$$4381/B2 sky130_fd_sc_hd__buf_4
Xrepeater686 U$$416/X VGND VGND VPWR VPWR U$$545/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_42_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater697 U$$4107/B2 VGND VGND VPWR VPWR U$$4081/B2 sky130_fd_sc_hd__buf_4
XFILLER_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4390 U$$4390/A1 U$$4388/X U$$4392/A1 U$$4389/X VGND VGND VPWR VPWR U$$4391/A sky130_fd_sc_hd__a22o_1
XFILLER_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_467 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_91_0 dadda_fa_4_91_0/A dadda_fa_4_91_0/B dadda_fa_4_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_92_0/A dadda_fa_5_91_1/A sky130_fd_sc_hd__fa_1
XFILLER_147_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_105_2 U$$4473/X input135/X dadda_fa_3_105_2/CIN VGND VGND VPWR VPWR dadda_fa_4_106_1/A
+ dadda_fa_4_105_2/B sky130_fd_sc_hd__fa_1
XFILLER_164_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_119_0 dadda_fa_6_119_0/A dadda_fa_6_119_0/B dadda_fa_6_119_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_120_0/B dadda_fa_7_119_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$800 U$$800/A U$$804/B VGND VGND VPWR VPWR U$$800/X sky130_fd_sc_hd__xor2_1
X_673_ _679_/CLK _673_/D VGND VGND VPWR VPWR _673_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$811 U$$811/A1 U$$819/A2 U$$950/A1 U$$819/B2 VGND VGND VPWR VPWR U$$812/A sky130_fd_sc_hd__a22o_1
XFILLER_90_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$822 _627_/Q VGND VGND VPWR VPWR U$$822/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_3_39_3 dadda_fa_3_39_3/A dadda_fa_3_39_3/B dadda_fa_3_39_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_1/B dadda_fa_4_39_2/CIN sky130_fd_sc_hd__fa_1
XU$$833 U$$833/A U$$859/B VGND VGND VPWR VPWR U$$833/X sky130_fd_sc_hd__xor2_1
XFILLER_21_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$844 U$$22/A1 U$$878/A2 U$$981/B1 U$$878/B2 VGND VGND VPWR VPWR U$$845/A sky130_fd_sc_hd__a22o_1
XU$$855 U$$855/A U$$925/B VGND VGND VPWR VPWR U$$855/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1005 U$$2375/A1 U$$979/A2 U$$48/A1 U$$979/B2 VGND VGND VPWR VPWR U$$1006/A sky130_fd_sc_hd__a22o_1
XU$$866 U$$866/A1 U$$896/A2 U$$866/B1 U$$896/B2 VGND VGND VPWR VPWR U$$867/A sky130_fd_sc_hd__a22o_1
XU$$877 U$$877/A U$$879/B VGND VGND VPWR VPWR U$$877/X sky130_fd_sc_hd__xor2_1
XFILLER_71_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1016 U$$1016/A U$$1040/B VGND VGND VPWR VPWR U$$1016/X sky130_fd_sc_hd__xor2_1
XFILLER_16_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$888 U$$66/A1 U$$928/A2 U$$66/B1 U$$928/B2 VGND VGND VPWR VPWR U$$889/A sky130_fd_sc_hd__a22o_1
XFILLER_44_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1027 U$$68/A1 U$$999/A2 U$$70/A1 U$$999/B2 VGND VGND VPWR VPWR U$$1028/A sky130_fd_sc_hd__a22o_1
XU$$1038 U$$1038/A U$$1040/B VGND VGND VPWR VPWR U$$1038/X sky130_fd_sc_hd__xor2_1
XU$$899 U$$899/A U$$907/B VGND VGND VPWR VPWR U$$899/X sky130_fd_sc_hd__xor2_1
XU$$1049 U$$912/A1 U$$1089/A2 U$$914/A1 U$$1089/B2 VGND VGND VPWR VPWR U$$1050/A sky130_fd_sc_hd__a22o_1
XFILLER_71_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1700 _553_/Q VGND VGND VPWR VPWR U$$556/B1 sky130_fd_sc_hd__buf_4
XFILLER_99_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_2_28_3 U$$1260/X U$$1393/X VGND VGND VPWR VPWR dadda_fa_3_29_2/CIN dadda_fa_4_28_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_6_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_41_3 U$$2749/X input192/X dadda_fa_2_41_3/CIN VGND VGND VPWR VPWR dadda_fa_3_42_1/B
+ dadda_fa_3_41_3/B sky130_fd_sc_hd__fa_1
XFILLER_19_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_304 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_34_2 U$$1139/X U$$1272/X U$$1405/X VGND VGND VPWR VPWR dadda_fa_3_35_1/A
+ dadda_fa_3_34_3/A sky130_fd_sc_hd__fa_1
XU$$2240 U$$2375/B1 U$$2242/A2 U$$3884/B1 U$$2242/B2 VGND VGND VPWR VPWR U$$2241/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_11_1 dadda_fa_5_11_1/A dadda_fa_5_11_1/B dadda_ha_4_11_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_12_0/B dadda_fa_7_11_0/A sky130_fd_sc_hd__fa_1
XFILLER_23_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2251 U$$2251/A U$$2303/B VGND VGND VPWR VPWR U$$2251/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_27_1 U$$460/X U$$593/X U$$726/X VGND VGND VPWR VPWR dadda_fa_3_28_2/B
+ dadda_fa_3_27_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2262 U$$890/B1 U$$2262/A2 U$$757/A1 U$$2262/B2 VGND VGND VPWR VPWR U$$2263/A sky130_fd_sc_hd__a22o_1
XFILLER_179_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2273 U$$2273/A U$$2309/B VGND VGND VPWR VPWR U$$2273/X sky130_fd_sc_hd__xor2_1
XFILLER_90_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2284 U$$914/A1 U$$2326/A2 U$$914/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2285/A sky130_fd_sc_hd__a22o_1
XFILLER_179_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2295 U$$2295/A U$$2299/B VGND VGND VPWR VPWR U$$2295/X sky130_fd_sc_hd__xor2_1
XU$$1550 U$$1550/A U$$1562/B VGND VGND VPWR VPWR U$$1550/X sky130_fd_sc_hd__xor2_1
XU$$1561 U$$52/B1 U$$1561/A2 U$$467/A1 U$$1561/B2 VGND VGND VPWR VPWR U$$1562/A sky130_fd_sc_hd__a22o_1
XU$$1572 U$$1572/A U$$1578/B VGND VGND VPWR VPWR U$$1572/X sky130_fd_sc_hd__xor2_1
XFILLER_72_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1583 U$$896/B1 U$$1587/A2 U$$900/A1 U$$1587/B2 VGND VGND VPWR VPWR U$$1584/A sky130_fd_sc_hd__a22o_1
XU$$1594 U$$1594/A U$$1598/B VGND VGND VPWR VPWR U$$1594/X sky130_fd_sc_hd__xor2_1
XFILLER_147_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_79_4 U$$2692/X U$$2825/X U$$2958/X VGND VGND VPWR VPWR dadda_fa_2_80_1/CIN
+ dadda_fa_2_79_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$202 final_adder.U$$697/A final_adder.U$$696/A VGND VGND VPWR VPWR
+ final_adder.U$$292/A sky130_fd_sc_hd__and2_1
XFILLER_131_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$213 final_adder.U$$707/A final_adder.U$$579/B1 final_adder.U$$213/B1
+ VGND VGND VPWR VPWR final_adder.U$$213/X sky130_fd_sc_hd__a21o_1
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$224 final_adder.U$$719/A final_adder.U$$718/A VGND VGND VPWR VPWR
+ final_adder.U$$304/B sky130_fd_sc_hd__and2_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_49_2 dadda_fa_4_49_2/A dadda_fa_4_49_2/B dadda_fa_4_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/CIN dadda_fa_5_49_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$235 final_adder.U$$729/A final_adder.U$$601/B1 final_adder.U$$235/B1
+ VGND VGND VPWR VPWR final_adder.U$$235/X sky130_fd_sc_hd__a21o_1
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$246 final_adder.U$$741/A final_adder.U$$740/A VGND VGND VPWR VPWR
+ final_adder.U$$314/A sky130_fd_sc_hd__and2_1
Xrepeater450 U$$4035/A2 VGND VGND VPWR VPWR U$$4005/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$257 final_adder.U$$130/X final_adder.U$$624/B final_adder.U$$131/X
+ VGND VGND VPWR VPWR final_adder.U$$626/B sky130_fd_sc_hd__a21o_1
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater461 U$$3840/X VGND VGND VPWR VPWR U$$3968/A2 sky130_fd_sc_hd__buf_6
XU$$107 U$$107/A U$$117/B VGND VGND VPWR VPWR U$$107/X sky130_fd_sc_hd__xor2_1
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater472 U$$3696/A2 VGND VGND VPWR VPWR U$$3636/A2 sky130_fd_sc_hd__buf_8
Xfinal_adder.U$$268 final_adder.U$$268/A final_adder.U$$268/B VGND VGND VPWR VPWR
+ final_adder.U$$326/B sky130_fd_sc_hd__and2_1
XFILLER_211_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$118 U$$253/B1 U$$118/A2 U$$942/A1 U$$118/B2 VGND VGND VPWR VPWR U$$119/A sky130_fd_sc_hd__a22o_1
XFILLER_45_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$279 final_adder.U$$278/A final_adder.U$$173/X final_adder.U$$175/X
+ VGND VGND VPWR VPWR final_adder.U$$279/X sky130_fd_sc_hd__a21o_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater483 U$$3545/A2 VGND VGND VPWR VPWR U$$3559/A2 sky130_fd_sc_hd__buf_4
XFILLER_84_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_19_0 dadda_fa_7_19_0/A dadda_fa_7_19_0/B dadda_fa_7_19_0/CIN VGND VGND
+ VPWR VPWR _444_/D _315_/D sky130_fd_sc_hd__fa_1
XU$$129 U$$129/A U$$129/B VGND VGND VPWR VPWR U$$129/X sky130_fd_sc_hd__xor2_1
Xrepeater494 U$$3285/A2 VGND VGND VPWR VPWR U$$3209/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_84_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1007 U$$2813/B VGND VGND VPWR VPWR U$$2787/B sky130_fd_sc_hd__buf_6
XFILLER_175_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_110_0 dadda_fa_3_110_0/A U$$3286/X U$$3419/X VGND VGND VPWR VPWR dadda_fa_4_111_0/CIN
+ dadda_fa_4_110_1/CIN sky130_fd_sc_hd__fa_1
Xrepeater1018 U$$2739/A VGND VGND VPWR VPWR U$$2734/B sky130_fd_sc_hd__buf_8
Xrepeater1029 U$$2462/B VGND VGND VPWR VPWR U$$2418/B sky130_fd_sc_hd__buf_6
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput220 c[67] VGND VGND VPWR VPWR input220/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput231 c[77] VGND VGND VPWR VPWR input231/X sky130_fd_sc_hd__buf_4
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_51_2 dadda_fa_3_51_2/A dadda_fa_3_51_2/B dadda_fa_3_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_1/A dadda_fa_4_51_2/B sky130_fd_sc_hd__fa_1
Xinput242 c[87] VGND VGND VPWR VPWR input242/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_67_2 U$$939/X U$$1072/X U$$1205/X VGND VGND VPWR VPWR dadda_fa_1_68_6/A
+ dadda_fa_1_67_8/A sky130_fd_sc_hd__fa_1
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput253 c[97] VGND VGND VPWR VPWR input253/X sky130_fd_sc_hd__clkbuf_4
XTAP_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_44_1 dadda_fa_3_44_1/A dadda_fa_3_44_1/B dadda_fa_3_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_0/CIN dadda_fa_4_44_2/A sky130_fd_sc_hd__fa_1
XTAP_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_21_0 dadda_fa_6_21_0/A dadda_fa_6_21_0/B dadda_fa_6_21_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_22_0/B dadda_fa_7_21_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_37_0 dadda_fa_3_37_0/A dadda_fa_3_37_0/B dadda_fa_3_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_0/B dadda_fa_4_37_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_656_ _660_/CLK _656_/D VGND VGND VPWR VPWR _656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$630 U$$82/A1 U$$632/A2 U$$84/A1 U$$632/B2 VGND VGND VPWR VPWR U$$631/A sky130_fd_sc_hd__a22o_1
XU$$641 U$$641/A U$$651/B VGND VGND VPWR VPWR U$$641/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$652 U$$924/B1 U$$682/A2 U$$791/A1 U$$682/B2 VGND VGND VPWR VPWR U$$653/A sky130_fd_sc_hd__a22o_1
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$663 U$$663/A U$$665/B VGND VGND VPWR VPWR U$$663/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$674 U$$674/A1 U$$552/X U$$950/A1 U$$553/X VGND VGND VPWR VPWR U$$675/A sky130_fd_sc_hd__a22o_1
X_587_ _596_/CLK _587_/D VGND VGND VPWR VPWR _587_/Q sky130_fd_sc_hd__dfxtp_2
XU$$685 U$$685/A VGND VGND VPWR VPWR U$$685/Y sky130_fd_sc_hd__inv_1
XFILLER_44_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$696 U$$696/A U$$726/B VGND VGND VPWR VPWR U$$696/X sky130_fd_sc_hd__xor2_1
XFILLER_16_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_96_4 U$$4056/X U$$4189/X U$$4322/X VGND VGND VPWR VPWR dadda_fa_3_97_1/CIN
+ dadda_fa_3_96_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1530 U$$4160/B1 VGND VGND VPWR VPWR U$$3475/B1 sky130_fd_sc_hd__buf_4
XFILLER_144_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1541 U$$4158/A1 VGND VGND VPWR VPWR U$$2375/B1 sky130_fd_sc_hd__buf_6
XFILLER_172_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1552 U$$4293/A1 VGND VGND VPWR VPWR U$$866/B1 sky130_fd_sc_hd__buf_4
XFILLER_158_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1563 _570_/Q VGND VGND VPWR VPWR U$$4154/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_89_3 input244/X dadda_fa_2_89_3/B dadda_fa_2_89_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_90_1/B dadda_fa_3_89_3/B sky130_fd_sc_hd__fa_1
Xrepeater1574 U$$451/A1 VGND VGND VPWR VPWR U$$999/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_113_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1585 U$$4285/A1 VGND VGND VPWR VPWR U$$2641/A1 sky130_fd_sc_hd__buf_4
XFILLER_119_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1596 U$$993/A1 VGND VGND VPWR VPWR U$$34/A1 sky130_fd_sc_hd__buf_6
XFILLER_141_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_919 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_59_1 dadda_fa_5_59_1/A dadda_fa_5_59_1/B dadda_fa_5_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_60_0/B dadda_fa_7_59_0/A sky130_fd_sc_hd__fa_2
XFILLER_101_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_105_1 U$$3276/X U$$3409/X U$$3542/X VGND VGND VPWR VPWR dadda_fa_3_106_3/B
+ dadda_fa_4_105_0/A sky130_fd_sc_hd__fa_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2070 U$$2070/A U$$2108/B VGND VGND VPWR VPWR U$$2070/X sky130_fd_sc_hd__xor2_1
XFILLER_126_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2081 U$$985/A1 U$$2145/A2 U$$987/A1 U$$2145/B2 VGND VGND VPWR VPWR U$$2082/A sky130_fd_sc_hd__a22o_1
XFILLER_211_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_392 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2092 U$$2092/A U$$2136/B VGND VGND VPWR VPWR U$$2092/X sky130_fd_sc_hd__xor2_1
XFILLER_11_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1380 U$$8/B1 U$$1428/A2 U$$12/A1 U$$1428/B2 VGND VGND VPWR VPWR U$$1381/A sky130_fd_sc_hd__a22o_1
XFILLER_210_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1391 U$$1391/A U$$1459/B VGND VGND VPWR VPWR U$$1391/X sky130_fd_sc_hd__xor2_1
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4459_1808 VGND VGND VPWR VPWR U$$4459_1808/HI U$$4459/B sky130_fd_sc_hd__conb_1
XFILLER_149_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_84_2 U$$2170/X U$$2303/X U$$2436/X VGND VGND VPWR VPWR dadda_fa_2_85_2/CIN
+ dadda_fa_2_84_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_61_1 dadda_fa_4_61_1/A dadda_fa_4_61_1/B dadda_fa_4_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/B dadda_fa_5_61_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_77_1 U$$1757/X U$$1890/X U$$2023/X VGND VGND VPWR VPWR dadda_fa_2_78_0/CIN
+ dadda_fa_2_77_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_54_0 dadda_fa_4_54_0/A dadda_fa_4_54_0/B dadda_fa_4_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/A dadda_fa_5_54_1/A sky130_fd_sc_hd__fa_1
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_510_ _510_/CLK _510_/D VGND VGND VPWR VPWR _510_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 _235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_314 _237_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_325 _238_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_336 U$$1095/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_441_ _441_/CLK _441_/D VGND VGND VPWR VPWR _441_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_347 U$$761/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_358 _619_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_369 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_372_ _372_/CLK _372_/D VGND VGND VPWR VPWR _372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_99_2 dadda_fa_3_99_2/A dadda_fa_3_99_2/B dadda_fa_3_99_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_1/A dadda_fa_4_99_2/B sky130_fd_sc_hd__fa_1
XFILLER_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_69_0 dadda_fa_6_69_0/A dadda_fa_6_69_0/B dadda_fa_6_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_70_0/B dadda_fa_7_69_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_72_0 dadda_fa_0_72_0/A U$$683/X U$$816/X VGND VGND VPWR VPWR dadda_fa_1_73_7/A
+ dadda_fa_1_72_8/A sky130_fd_sc_hd__fa_1
XFILLER_27_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$460 U$$460/A U$$532/B VGND VGND VPWR VPWR U$$460/X sky130_fd_sc_hd__xor2_1
X_639_ _642_/CLK _639_/D VGND VGND VPWR VPWR _639_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_51_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$471 U$$745/A1 U$$483/A2 U$$882/B1 U$$483/B2 VGND VGND VPWR VPWR U$$472/A sky130_fd_sc_hd__a22o_1
XU$$482 U$$482/A U$$484/B VGND VGND VPWR VPWR U$$482/X sky130_fd_sc_hd__xor2_1
XU$$493 U$$493/A1 U$$499/A2 U$$84/A1 U$$499/B2 VGND VGND VPWR VPWR U$$494/A sky130_fd_sc_hd__a22o_1
XFILLER_205_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_94_1 U$$3121/X U$$3254/X U$$3387/X VGND VGND VPWR VPWR dadda_fa_3_95_0/CIN
+ dadda_fa_3_94_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_71_0 dadda_fa_5_71_0/A dadda_fa_5_71_0/B dadda_fa_5_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_72_0/A dadda_fa_6_71_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1360 U$$3791/B1 VGND VGND VPWR VPWR U$$4065/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_87_0 U$$3639/X U$$3772/X U$$3905/X VGND VGND VPWR VPWR dadda_fa_3_88_0/B
+ dadda_fa_3_87_2/B sky130_fd_sc_hd__fa_1
Xrepeater1371 U$$2830/A1 VGND VGND VPWR VPWR U$$501/A1 sky130_fd_sc_hd__buf_6
XFILLER_158_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1382 U$$3650/A1 VGND VGND VPWR VPWR U$$2963/B1 sky130_fd_sc_hd__buf_8
Xrepeater1393 _591_/Q VGND VGND VPWR VPWR U$$4470/A1 sky130_fd_sc_hd__buf_6
XFILLER_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_70_8 dadda_fa_1_70_8/A dadda_fa_1_70_8/B dadda_fa_1_70_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_3/A dadda_fa_3_70_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_1_63_7 dadda_fa_1_63_7/A dadda_fa_1_63_7/B dadda_fa_1_63_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_2/CIN dadda_fa_2_63_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_56_6 U$$3577/X U$$3710/X U$$3843/X VGND VGND VPWR VPWR dadda_fa_2_57_2/B
+ dadda_fa_2_56_5/B sky130_fd_sc_hd__fa_1
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_49_5 U$$2100/X U$$2233/X U$$2366/X VGND VGND VPWR VPWR dadda_fa_2_50_2/B
+ dadda_fa_2_49_5/B sky130_fd_sc_hd__fa_1
XFILLER_131_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_8_0 dadda_fa_7_8_0/A dadda_fa_7_8_0/B dadda_fa_7_8_0/CIN VGND VGND VPWR
+ VPWR _433_/D _304_/D sky130_fd_sc_hd__fa_1
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_86_0 dadda_fa_7_86_0/A dadda_fa_7_86_0/B dadda_fa_7_86_0/CIN VGND VGND
+ VPWR VPWR _511_/D _382_/D sky130_fd_sc_hd__fa_1
XFILLER_137_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4513_1835 VGND VGND VPWR VPWR U$$4513_1835/HI U$$4513/B sky130_fd_sc_hd__conb_1
XFILLER_85_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1066 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4208 U$$4482/A1 U$$4114/X U$$4208/B1 U$$4115/X VGND VGND VPWR VPWR U$$4209/A sky130_fd_sc_hd__a22o_1
XFILLER_172_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4219 U$$4219/A U$$4246/A VGND VGND VPWR VPWR U$$4219/X sky130_fd_sc_hd__xor2_1
XFILLER_46_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3507 U$$3779/B1 U$$3429/X U$$3646/A1 U$$3430/X VGND VGND VPWR VPWR U$$3508/A sky130_fd_sc_hd__a22o_1
XFILLER_105_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3518 U$$3518/A U$$3520/B VGND VGND VPWR VPWR U$$3518/X sky130_fd_sc_hd__xor2_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_101_0 dadda_fa_6_101_0/A dadda_fa_6_101_0/B dadda_fa_6_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_102_0/B dadda_fa_7_101_0/CIN sky130_fd_sc_hd__fa_1
XU$$3529 U$$3529/A1 U$$3531/A2 U$$3805/A1 U$$3531/B2 VGND VGND VPWR VPWR U$$3530/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2806 U$$3902/A1 U$$2832/A2 U$$3902/B1 U$$2832/B2 VGND VGND VPWR VPWR U$$2807/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _287_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2817 U$$2817/A U$$2861/B VGND VGND VPWR VPWR U$$2817/X sky130_fd_sc_hd__xor2_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2828 U$$3650/A1 U$$2832/A2 U$$2830/A1 U$$2832/B2 VGND VGND VPWR VPWR U$$2829/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2839 U$$2839/A U$$2839/B VGND VGND VPWR VPWR U$$2839/X sky130_fd_sc_hd__xor2_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _290_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _180_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _183_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_424_ _442_/CLK _424_/D VGND VGND VPWR VPWR _424_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_177 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_188 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_199 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1056 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_355_ _484_/CLK _355_/D VGND VGND VPWR VPWR _355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_286_ _526_/CLK _286_/D VGND VGND VPWR VPWR _286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3431_1751 VGND VGND VPWR VPWR U$$3431_1751/HI U$$3431/A1 sky130_fd_sc_hd__conb_1
XFILLER_127_423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_66_5 dadda_fa_2_66_5/A dadda_fa_2_66_5/B dadda_fa_2_66_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_2/A dadda_fa_4_66_0/A sky130_fd_sc_hd__fa_1
XFILLER_116_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_59_4 dadda_fa_2_59_4/A dadda_fa_2_59_4/B dadda_fa_2_59_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/CIN dadda_fa_3_59_3/CIN sky130_fd_sc_hd__fa_1
XTAP_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 a[14] VGND VGND VPWR VPWR _630_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_49_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$290 U$$973/B1 U$$308/A2 U$$429/A1 U$$308/B2 VGND VGND VPWR VPWR U$$291/A sky130_fd_sc_hd__a22o_1
XFILLER_20_502 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$4 _428_/Q _300_/Q VGND VGND VPWR VPWR final_adder.U$$499/B1 final_adder.U$$626/A
+ sky130_fd_sc_hd__ha_1
XFILLER_195_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput310 _200_/Q VGND VGND VPWR VPWR o[32] sky130_fd_sc_hd__buf_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput321 _210_/Q VGND VGND VPWR VPWR o[42] sky130_fd_sc_hd__buf_2
XFILLER_156_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput332 _220_/Q VGND VGND VPWR VPWR o[52] sky130_fd_sc_hd__buf_2
XFILLER_195_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 _230_/Q VGND VGND VPWR VPWR o[62] sky130_fd_sc_hd__buf_2
Xoutput354 _240_/Q VGND VGND VPWR VPWR o[72] sky130_fd_sc_hd__buf_2
Xoutput365 _250_/Q VGND VGND VPWR VPWR o[82] sky130_fd_sc_hd__buf_2
Xoutput376 _260_/Q VGND VGND VPWR VPWR o[92] sky130_fd_sc_hd__buf_2
Xrepeater1190 U$$2/A VGND VGND VPWR VPWR U$$129/B sky130_fd_sc_hd__buf_6
XFILLER_102_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_4 U$$3587/X U$$3720/X U$$3853/X VGND VGND VPWR VPWR dadda_fa_2_62_1/CIN
+ dadda_fa_2_61_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_3 U$$1977/X U$$2110/X U$$2243/X VGND VGND VPWR VPWR dadda_fa_2_55_1/B
+ dadda_fa_2_54_4/B sky130_fd_sc_hd__fa_1
XFILLER_132_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_31_2 dadda_fa_4_31_2/A dadda_fa_4_31_2/B dadda_fa_4_31_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/CIN dadda_fa_5_31_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_47_2 U$$899/X U$$1032/X U$$1165/X VGND VGND VPWR VPWR dadda_fa_2_48_2/A
+ dadda_fa_2_47_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_24_1 dadda_fa_4_24_1/A dadda_fa_4_24_1/B dadda_fa_4_24_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/B dadda_fa_5_24_1/B sky130_fd_sc_hd__fa_1
XFILLER_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_17_0 U$$706/X U$$839/X U$$972/X VGND VGND VPWR VPWR dadda_fa_5_18_0/A
+ dadda_fa_5_17_1/A sky130_fd_sc_hd__fa_1
XFILLER_208_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3__f_clk clkbuf_2_1_0_clk/X VGND VGND VPWR VPWR _479_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_23 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_69_3 dadda_fa_3_69_3/A dadda_fa_3_69_3/B dadda_fa_3_69_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_1/B dadda_fa_4_69_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4005 U$$4140/B1 U$$4005/A2 U$$4007/A1 U$$4005/B2 VGND VGND VPWR VPWR U$$4006/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4016 U$$4016/A U$$4058/B VGND VGND VPWR VPWR U$$4016/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4027 U$$4027/A1 U$$4065/A2 U$$4027/B1 U$$4065/B2 VGND VGND VPWR VPWR U$$4028/A
+ sky130_fd_sc_hd__a22o_1
XU$$4038 U$$4038/A U$$4084/B VGND VGND VPWR VPWR U$$4038/X sky130_fd_sc_hd__xor2_1
XFILLER_93_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3304 U$$3578/A1 U$$3356/A2 U$$3578/B1 U$$3356/B2 VGND VGND VPWR VPWR U$$3305/A
+ sky130_fd_sc_hd__a22o_1
XU$$4049 U$$4186/A1 U$$4061/A2 U$$4051/A1 U$$4061/B2 VGND VGND VPWR VPWR U$$4050/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3315 U$$3315/A U$$3343/B VGND VGND VPWR VPWR U$$3315/X sky130_fd_sc_hd__xor2_1
XU$$3326 U$$3735/B1 U$$3368/A2 U$$3602/A1 U$$3368/B2 VGND VGND VPWR VPWR U$$3327/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3337 U$$3337/A U$$3424/A VGND VGND VPWR VPWR U$$3337/X sky130_fd_sc_hd__xor2_1
XFILLER_47_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2603 U$$2603/A VGND VGND VPWR VPWR U$$2603/Y sky130_fd_sc_hd__inv_1
XFILLER_202_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3348 U$$3485/A1 U$$3356/A2 U$$3624/A1 U$$3356/B2 VGND VGND VPWR VPWR U$$3349/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3359 U$$3359/A U$$3407/B VGND VGND VPWR VPWR U$$3359/X sky130_fd_sc_hd__xor2_1
XFILLER_47_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2614 U$$2614/A U$$2654/B VGND VGND VPWR VPWR U$$2614/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2625 U$$2625/A1 U$$2653/A2 U$$3584/B1 U$$2653/B2 VGND VGND VPWR VPWR U$$2626/A
+ sky130_fd_sc_hd__a22o_1
XU$$2636 U$$2636/A U$$2688/B VGND VGND VPWR VPWR U$$2636/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1902 U$$1902/A U$$1916/B VGND VGND VPWR VPWR U$$1902/X sky130_fd_sc_hd__xor2_1
XU$$2647 U$$3741/B1 U$$2653/A2 U$$4293/A1 U$$2653/B2 VGND VGND VPWR VPWR U$$2648/A
+ sky130_fd_sc_hd__a22o_1
XU$$2658 U$$2658/A U$$2664/B VGND VGND VPWR VPWR U$$2658/X sky130_fd_sc_hd__xor2_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1913 U$$2459/B1 U$$1915/A2 U$$545/A1 U$$1915/B2 VGND VGND VPWR VPWR U$$1914/A
+ sky130_fd_sc_hd__a22o_1
XU$$1924 U$$1924/A1 U$$1922/X U$$967/A1 U$$1923/X VGND VGND VPWR VPWR U$$1925/A sky130_fd_sc_hd__a22o_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2669 U$$3902/A1 U$$2705/A2 U$$3902/B1 U$$2705/B2 VGND VGND VPWR VPWR U$$2670/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1935 U$$1935/A U$$1977/B VGND VGND VPWR VPWR U$$1935/X sky130_fd_sc_hd__xor2_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1946 U$$848/B1 U$$2010/A2 U$$715/A1 U$$2010/B2 VGND VGND VPWR VPWR U$$1947/A sky130_fd_sc_hd__a22o_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1957 U$$1957/A U$$1957/B VGND VGND VPWR VPWR U$$1957/X sky130_fd_sc_hd__xor2_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1968 U$$50/A1 U$$1976/A2 U$$52/A1 U$$1976/B2 VGND VGND VPWR VPWR U$$1969/A sky130_fd_sc_hd__a22o_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ _628_/CLK _407_/D VGND VGND VPWR VPWR _407_/Q sky130_fd_sc_hd__dfxtp_1
XU$$1979 U$$1979/A U$$2029/B VGND VGND VPWR VPWR U$$1979/X sky130_fd_sc_hd__xor2_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_986 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_338_ _467_/CLK _338_/D VGND VGND VPWR VPWR _338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_269_ _520_/CLK _269_/D VGND VGND VPWR VPWR _269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_71_3 dadda_fa_2_71_3/A dadda_fa_2_71_3/B dadda_fa_2_71_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/B dadda_fa_3_71_3/B sky130_fd_sc_hd__fa_1
XFILLER_124_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_64_2 dadda_fa_2_64_2/A dadda_fa_2_64_2/B dadda_fa_2_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/A dadda_fa_3_64_3/A sky130_fd_sc_hd__fa_1
XFILLER_110_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater802 U$$2437/B2 VGND VGND VPWR VPWR U$$2395/B2 sky130_fd_sc_hd__buf_4
XFILLER_97_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$609 final_adder.U$$736/A final_adder.U$$736/B final_adder.U$$609/B1
+ VGND VGND VPWR VPWR final_adder.U$$737/B sky130_fd_sc_hd__a21o_1
XFILLER_42_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater813 U$$2318/B2 VGND VGND VPWR VPWR U$$2326/B2 sky130_fd_sc_hd__buf_4
XFILLER_84_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater824 U$$1982/B2 VGND VGND VPWR VPWR U$$1976/B2 sky130_fd_sc_hd__buf_4
XFILLER_38_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_41_1 dadda_fa_5_41_1/A dadda_fa_5_41_1/B dadda_fa_5_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_42_0/B dadda_fa_7_41_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_57_1 dadda_fa_2_57_1/A dadda_fa_2_57_1/B dadda_fa_2_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_0/CIN dadda_fa_3_57_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater835 U$$1915/B2 VGND VGND VPWR VPWR U$$1897/B2 sky130_fd_sc_hd__buf_6
XFILLER_99_1029 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater846 U$$1649/X VGND VGND VPWR VPWR U$$1778/B2 sky130_fd_sc_hd__buf_6
Xrepeater857 U$$263/B2 VGND VGND VPWR VPWR U$$219/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_5_34_0 dadda_fa_5_34_0/A dadda_fa_5_34_0/B dadda_fa_5_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_35_0/A dadda_fa_6_34_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater868 U$$1500/B2 VGND VGND VPWR VPWR U$$1486/B2 sky130_fd_sc_hd__buf_6
XU$$20 U$$20/A1 U$$8/A2 U$$20/B1 U$$8/B2 VGND VGND VPWR VPWR U$$21/A sky130_fd_sc_hd__a22o_1
XFILLER_37_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater879 U$$1238/X VGND VGND VPWR VPWR U$$1345/B2 sky130_fd_sc_hd__buf_6
XU$$31 U$$31/A U$$57/B VGND VGND VPWR VPWR U$$31/X sky130_fd_sc_hd__xor2_1
XU$$42 U$$42/A1 U$$68/A2 U$$42/B1 U$$68/B2 VGND VGND VPWR VPWR U$$43/A sky130_fd_sc_hd__a22o_1
XU$$53 U$$53/A U$$99/B VGND VGND VPWR VPWR U$$53/X sky130_fd_sc_hd__xor2_1
XU$$64 U$$64/A1 U$$4/X U$$66/A1 U$$5/X VGND VGND VPWR VPWR U$$65/A sky130_fd_sc_hd__a22o_1
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$75 U$$75/A U$$81/B VGND VGND VPWR VPWR U$$75/X sky130_fd_sc_hd__xor2_1
XU$$3860 _560_/Q U$$3970/A2 U$$4136/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3861/A sky130_fd_sc_hd__a22o_1
XFILLER_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3871 U$$3871/A U$$3873/B VGND VGND VPWR VPWR U$$3871/X sky130_fd_sc_hd__xor2_1
XFILLER_80_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3882 U$$4154/B1 U$$3916/A2 U$$4156/B1 U$$3916/B2 VGND VGND VPWR VPWR U$$3883/A
+ sky130_fd_sc_hd__a22o_1
XU$$86 U$$86/A1 U$$98/A2 U$$88/A1 U$$98/B2 VGND VGND VPWR VPWR U$$87/A sky130_fd_sc_hd__a22o_1
XFILLER_64_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$97 U$$97/A U$$99/B VGND VGND VPWR VPWR U$$97/X sky130_fd_sc_hd__xor2_1
XU$$3893 U$$3893/A U$$3933/B VGND VGND VPWR VPWR U$$3893/X sky130_fd_sc_hd__xor2_1
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_11 _178_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_22 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_33 _282_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_44 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_66 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_99 _287_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_79_2 dadda_fa_4_79_2/A dadda_fa_4_79_2/B dadda_fa_4_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/CIN dadda_fa_5_79_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_49_0 dadda_fa_7_49_0/A dadda_fa_7_49_0/B dadda_fa_7_49_0/CIN VGND VGND
+ VPWR VPWR _474_/D _345_/D sky130_fd_sc_hd__fa_2
XFILLER_43_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_52_0 U$$377/X U$$510/X U$$643/X VGND VGND VPWR VPWR dadda_fa_2_53_0/B
+ dadda_fa_2_52_3/B sky130_fd_sc_hd__fa_1
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1066 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1209 U$$1209/A U$$1209/B VGND VGND VPWR VPWR U$$1209/X sky130_fd_sc_hd__xor2_1
XFILLER_203_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_clk _369_/CLK VGND VGND VPWR VPWR _516_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_81_2 dadda_fa_3_81_2/A dadda_fa_3_81_2/B dadda_fa_3_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_1/A dadda_fa_4_81_2/B sky130_fd_sc_hd__fa_1
XFILLER_152_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_74_1 dadda_fa_3_74_1/A dadda_fa_3_74_1/B dadda_fa_3_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_0/CIN dadda_fa_4_74_2/A sky130_fd_sc_hd__fa_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_51_0 dadda_fa_6_51_0/A dadda_fa_6_51_0/B dadda_fa_6_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_52_0/B dadda_fa_7_51_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_67_0 dadda_fa_3_67_0/A dadda_fa_3_67_0/B dadda_fa_3_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_0/B dadda_fa_4_67_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3101 U$$3101/A U$$3145/B VGND VGND VPWR VPWR U$$3101/X sky130_fd_sc_hd__xor2_1
XFILLER_93_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3112 U$$3112/A1 U$$3132/A2 U$$3934/B1 U$$3132/B2 VGND VGND VPWR VPWR U$$3113/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_110_2 dadda_fa_4_110_2/A dadda_fa_4_110_2/B dadda_ha_3_110_3/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_111_0/CIN dadda_fa_5_110_1/CIN sky130_fd_sc_hd__fa_1
XU$$3123 U$$3123/A U$$3133/B VGND VGND VPWR VPWR U$$3123/X sky130_fd_sc_hd__xor2_1
XU$$3134 U$$3269/B1 U$$3144/A2 U$$3273/A1 U$$3144/B2 VGND VGND VPWR VPWR U$$3135/A
+ sky130_fd_sc_hd__a22o_1
XU$$2400 U$$2400/A U$$2400/B VGND VGND VPWR VPWR U$$2400/X sky130_fd_sc_hd__xor2_1
XFILLER_74_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3145 U$$3145/A U$$3145/B VGND VGND VPWR VPWR U$$3145/X sky130_fd_sc_hd__xor2_1
XU$$3156 U$$3154/B _661_/Q _662_/Q U$$3151/Y VGND VGND VPWR VPWR U$$3156/X sky130_fd_sc_hd__a22o_1
XU$$2411 U$$3096/A1 U$$2435/A2 U$$3096/B1 U$$2435/B2 VGND VGND VPWR VPWR U$$2412/A
+ sky130_fd_sc_hd__a22o_1
XU$$2422 U$$2422/A U$$2462/B VGND VGND VPWR VPWR U$$2422/X sky130_fd_sc_hd__xor2_1
XFILLER_74_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_103_1 dadda_fa_4_103_1/A dadda_fa_4_103_1/B dadda_fa_4_103_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/B dadda_fa_5_103_1/B sky130_fd_sc_hd__fa_1
XU$$3167 U$$3578/A1 U$$3215/A2 U$$3578/B1 U$$3215/B2 VGND VGND VPWR VPWR U$$3168/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3178 U$$3178/A U$$3232/B VGND VGND VPWR VPWR U$$3178/X sky130_fd_sc_hd__xor2_1
XFILLER_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2433 U$$924/B1 U$$2435/A2 U$$2435/A1 U$$2435/B2 VGND VGND VPWR VPWR U$$2434/A
+ sky130_fd_sc_hd__a22o_1
XU$$3189 U$$3735/B1 U$$3235/A2 U$$3602/A1 U$$3235/B2 VGND VGND VPWR VPWR U$$3190/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2444 U$$2444/A U$$2466/A VGND VGND VPWR VPWR U$$2444/X sky130_fd_sc_hd__xor2_1
XU$$1710 U$$3217/A1 U$$1710/A2 U$$3354/B1 U$$1710/B2 VGND VGND VPWR VPWR U$$1711/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2455 U$$948/A1 U$$2463/A2 _612_/Q U$$2463/B2 VGND VGND VPWR VPWR U$$2456/A sky130_fd_sc_hd__a22o_1
XU$$2466 U$$2466/A VGND VGND VPWR VPWR U$$2466/Y sky130_fd_sc_hd__inv_1
XU$$1721 U$$1721/A U$$1747/B VGND VGND VPWR VPWR U$$1721/X sky130_fd_sc_hd__xor2_1
XU$$1732 U$$88/A1 U$$1648/X U$$90/A1 U$$1649/X VGND VGND VPWR VPWR U$$1733/A sky130_fd_sc_hd__a22o_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2477 U$$2477/A U$$2517/B VGND VGND VPWR VPWR U$$2477/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1743 U$$1743/A U$$1773/B VGND VGND VPWR VPWR U$$1743/X sky130_fd_sc_hd__xor2_1
XU$$2488 U$$2625/A1 U$$2524/A2 U$$3584/B1 U$$2524/B2 VGND VGND VPWR VPWR U$$2489/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1754 U$$3124/A1 U$$1762/A2 U$$3124/B1 U$$1762/B2 VGND VGND VPWR VPWR U$$1755/A
+ sky130_fd_sc_hd__a22o_1
XU$$2499 U$$2499/A U$$2517/B VGND VGND VPWR VPWR U$$2499/X sky130_fd_sc_hd__xor2_1
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1765 U$$1765/A U$$1773/B VGND VGND VPWR VPWR U$$1765/X sky130_fd_sc_hd__xor2_1
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1776 U$$678/B1 U$$1778/A2 U$$4105/B1 U$$1778/B2 VGND VGND VPWR VPWR U$$1777/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1787 U$$1787/A1 U$$1859/A2 U$$2746/B1 U$$1859/B2 VGND VGND VPWR VPWR U$$1788/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_7_124_0 dadda_fa_7_124_0/A dadda_fa_7_124_0/B dadda_fa_7_124_0/CIN VGND
+ VGND VPWR VPWR _549_/D _420_/D sky130_fd_sc_hd__fa_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1798 U$$1798/A U$$1820/B VGND VGND VPWR VPWR U$$1798/X sky130_fd_sc_hd__xor2_1
XFILLER_203_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_clk _369_/CLK VGND VGND VPWR VPWR _500_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_187_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput20 a[27] VGND VGND VPWR VPWR _643_/D sky130_fd_sc_hd__clkbuf_1
Xinput31 a[37] VGND VGND VPWR VPWR _653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 a[47] VGND VGND VPWR VPWR _663_/D sky130_fd_sc_hd__clkbuf_1
Xinput53 a[57] VGND VGND VPWR VPWR _673_/D sky130_fd_sc_hd__clkbuf_1
Xinput64 a[9] VGND VGND VPWR VPWR _625_/D sky130_fd_sc_hd__clkbuf_2
Xinput75 b[19] VGND VGND VPWR VPWR _571_/D sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_5_89_1 dadda_fa_5_89_1/A dadda_fa_5_89_1/B dadda_fa_5_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_90_0/B dadda_fa_7_89_0/A sky130_fd_sc_hd__fa_1
XFILLER_122_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput86 b[29] VGND VGND VPWR VPWR _581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput97 b[39] VGND VGND VPWR VPWR _591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater610 U$$263/A2 VGND VGND VPWR VPWR U$$195/A2 sky130_fd_sc_hd__buf_2
XFILLER_111_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$417 final_adder.U$$334/B final_adder.U$$678/B final_adder.U$$285/X
+ VGND VGND VPWR VPWR final_adder.U$$682/B sky130_fd_sc_hd__a21o_1
Xrepeater621 U$$1478/A2 VGND VGND VPWR VPWR U$$1500/A2 sky130_fd_sc_hd__buf_8
XFILLER_111_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater632 U$$1190/A2 VGND VGND VPWR VPWR U$$1150/A2 sky130_fd_sc_hd__buf_6
Xrepeater643 U$$997/B2 VGND VGND VPWR VPWR U$$999/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$439 final_adder.U$$262/B final_adder.U$$634/B final_adder.U$$141/X
+ VGND VGND VPWR VPWR final_adder.U$$636/B sky130_fd_sc_hd__a21o_1
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater654 U$$948/B2 VGND VGND VPWR VPWR U$$956/B2 sky130_fd_sc_hd__buf_6
Xrepeater665 U$$632/B2 VGND VGND VPWR VPWR U$$616/B2 sky130_fd_sc_hd__buf_4
Xrepeater676 U$$4345/B2 VGND VGND VPWR VPWR U$$4347/B2 sky130_fd_sc_hd__buf_4
Xrepeater687 U$$4174/B2 VGND VGND VPWR VPWR U$$4140/B2 sky130_fd_sc_hd__buf_4
XU$$4380 U$$4380/A U$$4382/B VGND VGND VPWR VPWR U$$4380/X sky130_fd_sc_hd__xor2_1
Xrepeater698 U$$3978/X VGND VGND VPWR VPWR U$$4107/B2 sky130_fd_sc_hd__buf_4
XU$$4391 U$$4391/A U$$4391/B VGND VGND VPWR VPWR U$$4391/X sky130_fd_sc_hd__xor2_1
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3690 U$$4238/A1 U$$3696/A2 U$$4238/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3691/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_1119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_91_1 dadda_fa_4_91_1/A dadda_fa_4_91_1/B dadda_fa_4_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_92_0/B dadda_fa_5_91_1/B sky130_fd_sc_hd__fa_1
XFILLER_193_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_84_0 dadda_fa_4_84_0/A dadda_fa_4_84_0/B dadda_fa_4_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/A dadda_fa_5_84_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_105_3 dadda_fa_3_105_3/A dadda_fa_3_105_3/B dadda_fa_3_105_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_106_1/B dadda_fa_4_105_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_clk _634_/CLK VGND VGND VPWR VPWR _496_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_672_ _679_/CLK _672_/D VGND VGND VPWR VPWR _672_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$801 U$$938/A1 U$$689/X U$$938/B1 U$$690/X VGND VGND VPWR VPWR U$$802/A sky130_fd_sc_hd__a22o_1
XFILLER_91_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$812 U$$812/A U$$821/A VGND VGND VPWR VPWR U$$812/X sky130_fd_sc_hd__xor2_1
XTAP_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$823 _628_/Q VGND VGND VPWR VPWR U$$825/B sky130_fd_sc_hd__inv_1
XFILLER_112_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$834 U$$971/A1 U$$860/A2 U$$973/A1 U$$860/B2 VGND VGND VPWR VPWR U$$835/A sky130_fd_sc_hd__a22o_1
Xdadda_ha_4_122_0_1877 VGND VGND VPWR VPWR dadda_ha_4_122_0/A dadda_ha_4_122_0_1877/LO
+ sky130_fd_sc_hd__conb_1
XU$$845 U$$845/A U$$879/B VGND VGND VPWR VPWR U$$845/X sky130_fd_sc_hd__xor2_1
XU$$856 U$$34/A1 U$$928/A2 U$$856/B1 U$$928/B2 VGND VGND VPWR VPWR U$$857/A sky130_fd_sc_hd__a22o_1
XFILLER_189_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1006 U$$1006/A U$$980/B VGND VGND VPWR VPWR U$$1006/X sky130_fd_sc_hd__xor2_1
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$867 U$$867/A U$$897/B VGND VGND VPWR VPWR U$$867/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1017 U$$58/A1 U$$1065/A2 U$$60/A1 U$$1065/B2 VGND VGND VPWR VPWR U$$1018/A sky130_fd_sc_hd__a22o_1
XU$$878 U$$878/A1 U$$878/A2 U$$880/A1 U$$878/B2 VGND VGND VPWR VPWR U$$879/A sky130_fd_sc_hd__a22o_1
XU$$889 U$$889/A U$$929/B VGND VGND VPWR VPWR U$$889/X sky130_fd_sc_hd__xor2_1
XU$$1028 U$$1028/A U$$982/B VGND VGND VPWR VPWR U$$1028/X sky130_fd_sc_hd__xor2_1
XFILLER_189_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1039 U$$80/A1 U$$1039/A2 U$$80/B1 U$$1039/B2 VGND VGND VPWR VPWR U$$1040/A sky130_fd_sc_hd__a22o_1
XFILLER_73_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk _432_/CLK VGND VGND VPWR VPWR _179_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_99_0 dadda_fa_6_99_0/A dadda_fa_6_99_0/B dadda_fa_6_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_100_0/B dadda_fa_7_99_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_156_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1701 _553_/Q VGND VGND VPWR VPWR U$$3709/A1 sky130_fd_sc_hd__buf_6
XFILLER_153_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_41_4 dadda_fa_2_41_4/A dadda_fa_2_41_4/B dadda_fa_2_41_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_42_1/CIN dadda_fa_3_41_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_208_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_34_3 U$$1538/X U$$1671/X U$$1804/X VGND VGND VPWR VPWR dadda_fa_3_35_1/B
+ dadda_fa_3_34_3/B sky130_fd_sc_hd__fa_1
XFILLER_34_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2230 U$$449/A1 U$$2248/A2 U$$449/B1 U$$2248/B2 VGND VGND VPWR VPWR U$$2231/A sky130_fd_sc_hd__a22o_1
XFILLER_34_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2241 U$$2241/A U$$2241/B VGND VGND VPWR VPWR U$$2241/X sky130_fd_sc_hd__xor2_1
XU$$2252 U$$4031/B1 U$$2302/A2 U$$3896/B1 U$$2302/B2 VGND VGND VPWR VPWR U$$2253/A
+ sky130_fd_sc_hd__a22o_1
XU$$2263 U$$2263/A U$$2263/B VGND VGND VPWR VPWR U$$2263/X sky130_fd_sc_hd__xor2_1
XFILLER_22_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2274 U$$3096/A1 U$$2274/A2 U$$3372/A1 U$$2274/B2 VGND VGND VPWR VPWR U$$2275/A
+ sky130_fd_sc_hd__a22o_1
XU$$1540 U$$1540/A U$$1578/B VGND VGND VPWR VPWR U$$1540/X sky130_fd_sc_hd__xor2_1
XU$$2285 U$$2285/A U$$2328/A VGND VGND VPWR VPWR U$$2285/X sky130_fd_sc_hd__xor2_1
XFILLER_179_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2296 U$$3529/A1 U$$2318/A2 U$$2435/A1 U$$2318/B2 VGND VGND VPWR VPWR U$$2297/A
+ sky130_fd_sc_hd__a22o_1
XU$$1551 U$$42/B1 U$$1557/A2 U$$729/B1 U$$1557/B2 VGND VGND VPWR VPWR U$$1552/A sky130_fd_sc_hd__a22o_1
XFILLER_179_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1562 U$$1562/A U$$1562/B VGND VGND VPWR VPWR U$$1562/X sky130_fd_sc_hd__xor2_1
XFILLER_195_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1573 U$$3217/A1 U$$1577/A2 U$$3354/B1 U$$1577/B2 VGND VGND VPWR VPWR U$$1574/A
+ sky130_fd_sc_hd__a22o_1
XU$$1584 U$$1584/A U$$1588/B VGND VGND VPWR VPWR U$$1584/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_14_clk _616_/CLK VGND VGND VPWR VPWR _343_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1595 U$$88/A1 U$$1597/A2 U$$90/A1 U$$1597/B2 VGND VGND VPWR VPWR U$$1596/A sky130_fd_sc_hd__a22o_1
XFILLER_176_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_955 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1008 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_79_5 U$$3091/X U$$3224/X U$$3357/X VGND VGND VPWR VPWR dadda_fa_2_80_2/A
+ dadda_fa_2_79_5/A sky130_fd_sc_hd__fa_1
XFILLER_44_1112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$203 final_adder.U$$697/A final_adder.U$$569/B1 final_adder.U$$203/B1
+ VGND VGND VPWR VPWR final_adder.U$$203/X sky130_fd_sc_hd__a21o_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$214 final_adder.U$$709/A final_adder.U$$708/A VGND VGND VPWR VPWR
+ final_adder.U$$298/A sky130_fd_sc_hd__and2_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$225 final_adder.U$$719/A final_adder.U$$591/B1 final_adder.U$$225/B1
+ VGND VGND VPWR VPWR final_adder.U$$225/X sky130_fd_sc_hd__a21o_1
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater440 U$$68/A2 VGND VGND VPWR VPWR U$$52/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$236 final_adder.U$$731/A final_adder.U$$730/A VGND VGND VPWR VPWR
+ final_adder.U$$310/B sky130_fd_sc_hd__and2_1
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$247 final_adder.U$$741/A final_adder.U$$613/B1 final_adder.U$$247/B1
+ VGND VGND VPWR VPWR final_adder.U$$247/X sky130_fd_sc_hd__a21o_1
Xrepeater451 U$$4095/A2 VGND VGND VPWR VPWR U$$4035/A2 sky130_fd_sc_hd__buf_6
XFILLER_100_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$258 final_adder.U$$258/A final_adder.U$$258/B VGND VGND VPWR VPWR
+ final_adder.U$$258/X sky130_fd_sc_hd__and2_1
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater462 U$$3769/A2 VGND VGND VPWR VPWR U$$3743/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$108 U$$517/B1 U$$118/A2 U$$382/B1 U$$118/B2 VGND VGND VPWR VPWR U$$109/A sky130_fd_sc_hd__a22o_1
Xrepeater473 U$$3688/A2 VGND VGND VPWR VPWR U$$3696/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$269 final_adder.U$$268/A final_adder.U$$153/X final_adder.U$$155/X
+ VGND VGND VPWR VPWR final_adder.U$$269/X sky130_fd_sc_hd__a21o_1
XU$$119 U$$119/A U$$129/B VGND VGND VPWR VPWR U$$119/X sky130_fd_sc_hd__xor2_1
Xrepeater484 U$$3555/A2 VGND VGND VPWR VPWR U$$3545/A2 sky130_fd_sc_hd__buf_4
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater495 U$$3285/A2 VGND VGND VPWR VPWR U$$3235/A2 sky130_fd_sc_hd__buf_6
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_616 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4401_1779 VGND VGND VPWR VPWR U$$4401_1779/HI U$$4401/B sky130_fd_sc_hd__conb_1
XFILLER_166_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_110_1 U$$3552/X U$$3685/X U$$3818/X VGND VGND VPWR VPWR dadda_fa_4_111_1/A
+ dadda_fa_4_110_2/A sky130_fd_sc_hd__fa_1
Xrepeater1008 U$$2843/B VGND VGND VPWR VPWR U$$2813/B sky130_fd_sc_hd__buf_8
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1019 U$$2739/A VGND VGND VPWR VPWR U$$2708/B sky130_fd_sc_hd__buf_12
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_103_0 U$$3937/X U$$4070/X U$$4203/X VGND VGND VPWR VPWR dadda_fa_4_104_0/B
+ dadda_fa_4_103_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_68_5 U$$2271/X U$$2404/X VGND VGND VPWR VPWR dadda_fa_1_69_7/B dadda_fa_2_68_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_108_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput210 c[58] VGND VGND VPWR VPWR input210/X sky130_fd_sc_hd__buf_2
XFILLER_88_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput221 c[68] VGND VGND VPWR VPWR input221/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput232 c[78] VGND VGND VPWR VPWR input232/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_51_3 dadda_fa_3_51_3/A dadda_fa_3_51_3/B dadda_fa_3_51_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_1/B dadda_fa_4_51_2/CIN sky130_fd_sc_hd__fa_1
Xinput243 c[88] VGND VGND VPWR VPWR input243/X sky130_fd_sc_hd__clkbuf_2
XTAP_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_67_3 U$$1338/X U$$1471/X U$$1604/X VGND VGND VPWR VPWR dadda_fa_1_68_6/B
+ dadda_fa_1_67_8/B sky130_fd_sc_hd__fa_1
Xinput254 c[98] VGND VGND VPWR VPWR input254/X sky130_fd_sc_hd__buf_4
XTAP_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_44_2 dadda_fa_3_44_2/A dadda_fa_3_44_2/B dadda_fa_3_44_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_1/A dadda_fa_4_44_2/B sky130_fd_sc_hd__fa_1
XFILLER_208_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_37_1 dadda_fa_3_37_1/A dadda_fa_3_37_1/B dadda_fa_3_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_0/CIN dadda_fa_4_37_2/A sky130_fd_sc_hd__fa_1
XU$$620 U$$757/A1 U$$668/A2 U$$759/A1 U$$670/B2 VGND VGND VPWR VPWR U$$621/A sky130_fd_sc_hd__a22o_1
XFILLER_84_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_655_ _662_/CLK _655_/D VGND VGND VPWR VPWR _655_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$631 U$$631/A U$$659/B VGND VGND VPWR VPWR U$$631/X sky130_fd_sc_hd__xor2_1
XU$$642 U$$914/B1 U$$650/A2 U$$916/B1 U$$650/B2 VGND VGND VPWR VPWR U$$643/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_14_0 dadda_fa_6_14_0/A dadda_fa_6_14_0/B dadda_fa_6_14_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_15_0/B dadda_fa_7_14_0/CIN sky130_fd_sc_hd__fa_1
XU$$653 U$$653/A U$$684/A VGND VGND VPWR VPWR U$$653/X sky130_fd_sc_hd__xor2_1
XFILLER_186_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1069 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$664 U$$938/A1 U$$668/A2 U$$938/B1 U$$670/B2 VGND VGND VPWR VPWR U$$665/A sky130_fd_sc_hd__a22o_1
XFILLER_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$675 U$$675/A U$$685/A VGND VGND VPWR VPWR U$$675/X sky130_fd_sc_hd__xor2_1
XFILLER_189_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_586_ _588_/CLK _586_/D VGND VGND VPWR VPWR _586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$686 _626_/Q VGND VGND VPWR VPWR U$$688/B sky130_fd_sc_hd__inv_1
XFILLER_210_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$697 U$$971/A1 U$$725/A2 U$$973/A1 U$$725/B2 VGND VGND VPWR VPWR U$$698/A sky130_fd_sc_hd__a22o_1
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_96_5 U$$4455/X input252/X dadda_fa_2_96_5/CIN VGND VGND VPWR VPWR dadda_fa_3_97_2/A
+ dadda_fa_4_96_0/A sky130_fd_sc_hd__fa_2
Xrepeater1520 U$$54/A1 VGND VGND VPWR VPWR U$$463/B1 sky130_fd_sc_hd__buf_4
Xrepeater1531 _574_/Q VGND VGND VPWR VPWR U$$4160/B1 sky130_fd_sc_hd__buf_4
XFILLER_158_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1542 U$$2786/B1 VGND VGND VPWR VPWR U$$733/A1 sky130_fd_sc_hd__buf_6
XFILLER_181_980 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1553 U$$4293/A1 VGND VGND VPWR VPWR U$$4430/A1 sky130_fd_sc_hd__buf_6
XFILLER_193_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_89_4 dadda_fa_2_89_4/A dadda_fa_2_89_4/B dadda_fa_2_89_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_90_1/CIN dadda_fa_3_89_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1564 U$$999/B1 VGND VGND VPWR VPWR U$$316/A1 sky130_fd_sc_hd__buf_8
XFILLER_158_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1575 U$$4287/A1 VGND VGND VPWR VPWR U$$451/A1 sky130_fd_sc_hd__buf_6
XFILLER_113_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1586 _567_/Q VGND VGND VPWR VPWR U$$4285/A1 sky130_fd_sc_hd__buf_6
XFILLER_99_747 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1597 U$$3320/B1 VGND VGND VPWR VPWR U$$993/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_67_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_clk _442_/CLK VGND VGND VPWR VPWR _454_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_32_0 U$$71/X U$$204/X U$$337/X VGND VGND VPWR VPWR dadda_fa_3_33_0/B dadda_fa_3_32_2/B
+ sky130_fd_sc_hd__fa_1
XFILLER_207_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2060 U$$2058/B _645_/Q _646_/Q U$$2055/Y VGND VGND VPWR VPWR U$$2060/X sky130_fd_sc_hd__a22o_4
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2071 U$$2345/A1 U$$2109/A2 U$$2895/A1 U$$2109/B2 VGND VGND VPWR VPWR U$$2072/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2082 U$$2082/A U$$2144/B VGND VGND VPWR VPWR U$$2082/X sky130_fd_sc_hd__xor2_1
XFILLER_195_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2093 U$$3187/B1 U$$2145/A2 U$$999/A1 U$$2145/B2 VGND VGND VPWR VPWR U$$2094/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_161_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1370 U$$1370/A VGND VGND VPWR VPWR U$$1370/Y sky130_fd_sc_hd__inv_1
XU$$1381 U$$1381/A U$$1429/B VGND VGND VPWR VPWR U$$1381/X sky130_fd_sc_hd__xor2_1
XU$$1392 U$$568/B1 U$$1458/A2 U$$435/A1 U$$1458/B2 VGND VGND VPWR VPWR U$$1393/A sky130_fd_sc_hd__a22o_1
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_119_0 input150/X dadda_fa_5_119_0/B dadda_fa_5_119_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_6_120_0/A dadda_fa_6_119_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_164_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_84_3 U$$2569/X U$$2702/X U$$2835/X VGND VGND VPWR VPWR dadda_fa_2_85_3/A
+ dadda_fa_2_84_5/A sky130_fd_sc_hd__fa_1
XFILLER_143_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_61_2 dadda_fa_4_61_2/A dadda_fa_4_61_2/B dadda_fa_4_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/CIN dadda_fa_5_61_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_77_2 U$$2156/X U$$2289/X U$$2422/X VGND VGND VPWR VPWR dadda_fa_2_78_1/A
+ dadda_fa_2_77_4/A sky130_fd_sc_hd__fa_1
XFILLER_98_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_54_1 dadda_fa_4_54_1/A dadda_fa_4_54_1/B dadda_fa_4_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/B dadda_fa_5_54_1/B sky130_fd_sc_hd__fa_1
XFILLER_98_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_730 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_31_0 dadda_fa_7_31_0/A dadda_fa_7_31_0/B dadda_fa_7_31_0/CIN VGND VGND
+ VPWR VPWR _456_/D _327_/D sky130_fd_sc_hd__fa_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_47_0 dadda_fa_4_47_0/A dadda_fa_4_47_0/B dadda_fa_4_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/A dadda_fa_5_47_1/A sky130_fd_sc_hd__fa_1
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_474 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_304 _235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_315 _237_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 _238_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_440_ _441_/CLK _440_/D VGND VGND VPWR VPWR _440_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_337 _560_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_348 U$$3503/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_359 U$$924/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_371_ _500_/CLK _371_/D VGND VGND VPWR VPWR _371_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_590 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4399_1778 VGND VGND VPWR VPWR U$$4399_1778/HI U$$4399/B sky130_fd_sc_hd__conb_1
XFILLER_210_892 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_99_3 dadda_fa_3_99_3/A dadda_fa_3_99_3/B dadda_fa_3_99_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_1/B dadda_fa_4_99_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_182_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_72_1 U$$949/X U$$1082/X U$$1215/X VGND VGND VPWR VPWR dadda_fa_1_73_7/B
+ dadda_fa_1_72_8/B sky130_fd_sc_hd__fa_1
XFILLER_209_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_65_0 _617_/Q U$$270/X U$$403/X VGND VGND VPWR VPWR dadda_fa_1_66_5/B dadda_fa_1_65_7/B
+ sky130_fd_sc_hd__fa_1
XFILLER_97_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$450 U$$450/A U$$484/B VGND VGND VPWR VPWR U$$450/X sky130_fd_sc_hd__xor2_1
X_638_ _642_/CLK _638_/D VGND VGND VPWR VPWR _638_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$461 U$$596/B1 U$$491/A2 U$$463/A1 U$$491/B2 VGND VGND VPWR VPWR U$$462/A sky130_fd_sc_hd__a22o_1
XFILLER_205_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$472 U$$472/A U$$484/B VGND VGND VPWR VPWR U$$472/X sky130_fd_sc_hd__xor2_1
XU$$483 U$$894/A1 U$$483/A2 U$$896/A1 U$$483/B2 VGND VGND VPWR VPWR U$$484/A sky130_fd_sc_hd__a22o_1
XFILLER_204_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$494 U$$494/A U$$500/B VGND VGND VPWR VPWR U$$494/X sky130_fd_sc_hd__xor2_1
XFILLER_32_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_569_ _569_/CLK _569_/D VGND VGND VPWR VPWR _569_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4423_1790 VGND VGND VPWR VPWR U$$4423_1790/HI U$$4423/B sky130_fd_sc_hd__conb_1
XFILLER_118_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_94_2 U$$3520/X U$$3653/X U$$3786/X VGND VGND VPWR VPWR dadda_fa_3_95_1/A
+ dadda_fa_3_94_3/A sky130_fd_sc_hd__fa_1
XFILLER_201_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_71_1 dadda_fa_5_71_1/A dadda_fa_5_71_1/B dadda_fa_5_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_72_0/B dadda_fa_7_71_0/A sky130_fd_sc_hd__fa_1
Xrepeater1350 U$$3932/A1 VGND VGND VPWR VPWR U$$3245/B1 sky130_fd_sc_hd__buf_6
Xrepeater1361 _595_/Q VGND VGND VPWR VPWR U$$4478/A1 sky130_fd_sc_hd__buf_4
XFILLER_114_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_87_1 U$$4038/X U$$4171/X U$$4304/X VGND VGND VPWR VPWR dadda_fa_3_88_0/CIN
+ dadda_fa_3_87_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_119_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1372 U$$3652/A1 VGND VGND VPWR VPWR U$$2830/A1 sky130_fd_sc_hd__buf_6
XFILLER_114_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1383 U$$4061/A1 VGND VGND VPWR VPWR U$$3650/A1 sky130_fd_sc_hd__buf_6
XFILLER_113_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1394 _591_/Q VGND VGND VPWR VPWR U$$4194/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_64_0 dadda_fa_5_64_0/A dadda_fa_5_64_0/B dadda_fa_5_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_65_0/A dadda_fa_6_64_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_119_1043 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_899 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_63_8 dadda_fa_1_63_8/A dadda_fa_1_63_8/B dadda_fa_1_63_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_3/A dadda_fa_3_63_0/A sky130_fd_sc_hd__fa_2
XFILLER_45_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_56_7 U$$3895/B input208/X dadda_fa_1_56_7/CIN VGND VGND VPWR VPWR dadda_fa_2_57_2/CIN
+ dadda_fa_2_56_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_49_6 U$$2499/X U$$2632/X U$$2765/X VGND VGND VPWR VPWR dadda_fa_2_50_2/CIN
+ dadda_fa_2_49_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_209_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_606 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_1_90_3 U$$2980/X U$$3113/X VGND VGND VPWR VPWR dadda_fa_2_91_5/A dadda_fa_3_90_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_148_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_79_0 dadda_fa_7_79_0/A dadda_fa_7_79_0/B dadda_fa_7_79_0/CIN VGND VGND
+ VPWR VPWR _504_/D _375_/D sky130_fd_sc_hd__fa_1
XFILLER_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_47 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_416 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_82_0 dadda_fa_1_82_0/A U$$1368/X U$$1501/X VGND VGND VPWR VPWR dadda_fa_2_83_1/B
+ dadda_fa_2_82_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_85_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4209 U$$4209/A U$$4215/B VGND VGND VPWR VPWR U$$4209/X sky130_fd_sc_hd__xor2_1
XFILLER_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3508 U$$3508/A U$$3562/A VGND VGND VPWR VPWR U$$3508/X sky130_fd_sc_hd__xor2_1
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3519 U$$916/A1 U$$3519/A2 U$$3519/B1 U$$3519/B2 VGND VGND VPWR VPWR U$$3520/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2807 U$$2807/A U$$2839/B VGND VGND VPWR VPWR U$$2807/X sky130_fd_sc_hd__xor2_1
XFILLER_73_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _287_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2818 U$$4051/A1 U$$2856/A2 U$$2957/A1 U$$2856/B2 VGND VGND VPWR VPWR U$$2819/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_455 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2829 U$$2829/A U$$2843/B VGND VGND VPWR VPWR U$$2829/X sky130_fd_sc_hd__xor2_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _290_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _180_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_423_ _550_/CLK _423_/D VGND VGND VPWR VPWR _423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_167 _183_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_178 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_354_ _484_/CLK _354_/D VGND VGND VPWR VPWR _354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_285_ _526_/CLK _285_/D VGND VGND VPWR VPWR _285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_81_0 dadda_fa_6_81_0/A dadda_fa_6_81_0/B dadda_fa_6_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_82_0/B dadda_fa_7_81_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_97_0 dadda_fa_3_97_0/A dadda_fa_3_97_0/B dadda_fa_3_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_0/B dadda_fa_4_97_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_182_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_858 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1031 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_59_5 dadda_fa_2_59_5/A dadda_fa_2_59_5/B dadda_fa_2_59_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_2/A dadda_fa_4_59_0/A sky130_fd_sc_hd__fa_2
XTAP_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 a[15] VGND VGND VPWR VPWR _631_/D sky130_fd_sc_hd__clkbuf_2
XTAP_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_731 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$280 U$$280/A1 U$$318/A2 U$$8/A1 U$$318/B2 VGND VGND VPWR VPWR U$$281/A sky130_fd_sc_hd__a22o_1
XFILLER_45_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$291 U$$291/A U$$309/B VGND VGND VPWR VPWR U$$291/X sky130_fd_sc_hd__xor2_1
XFILLER_178_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$5 _429_/Q _301_/Q VGND VGND VPWR VPWR final_adder.U$$5/COUT final_adder.U$$627/A
+ sky130_fd_sc_hd__ha_1
XFILLER_146_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput300 _191_/Q VGND VGND VPWR VPWR o[23] sky130_fd_sc_hd__buf_2
XFILLER_195_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput311 _201_/Q VGND VGND VPWR VPWR o[33] sky130_fd_sc_hd__buf_2
XFILLER_160_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput322 _211_/Q VGND VGND VPWR VPWR o[43] sky130_fd_sc_hd__buf_2
XFILLER_156_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput333 _221_/Q VGND VGND VPWR VPWR o[53] sky130_fd_sc_hd__buf_2
Xoutput344 _231_/Q VGND VGND VPWR VPWR o[63] sky130_fd_sc_hd__buf_2
XFILLER_195_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput355 _241_/Q VGND VGND VPWR VPWR o[73] sky130_fd_sc_hd__buf_2
Xrepeater1180 U$$272/B VGND VGND VPWR VPWR U$$264/B sky130_fd_sc_hd__buf_6
Xoutput366 _251_/Q VGND VGND VPWR VPWR o[83] sky130_fd_sc_hd__buf_2
Xoutput377 _261_/Q VGND VGND VPWR VPWR o[93] sky130_fd_sc_hd__buf_2
Xrepeater1191 _617_/Q VGND VGND VPWR VPWR U$$2/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_5 U$$3986/X U$$4119/X input214/X VGND VGND VPWR VPWR dadda_fa_2_62_2/A
+ dadda_fa_2_61_5/A sky130_fd_sc_hd__fa_1
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_54_4 U$$2376/X U$$2509/X U$$2642/X VGND VGND VPWR VPWR dadda_fa_2_55_1/CIN
+ dadda_fa_2_54_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_47_3 U$$1298/X U$$1431/X U$$1564/X VGND VGND VPWR VPWR dadda_fa_2_48_2/B
+ dadda_fa_2_47_5/A sky130_fd_sc_hd__fa_1
XFILLER_43_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_24_2 dadda_fa_4_24_2/A dadda_fa_4_24_2/B dadda_fa_4_24_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/CIN dadda_fa_5_24_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_17_1 U$$1105/X input165/X dadda_fa_4_17_1/CIN VGND VGND VPWR VPWR dadda_fa_5_18_0/B
+ dadda_fa_5_17_1/B sky130_fd_sc_hd__fa_1
XFILLER_24_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_1019 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_23 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_3_20_3 U$$1244/X U$$1377/X VGND VGND VPWR VPWR dadda_fa_4_21_1/B dadda_ha_3_20_3/SUM
+ sky130_fd_sc_hd__ha_1
XU$$4006 U$$4006/A U$$4036/B VGND VGND VPWR VPWR U$$4006/X sky130_fd_sc_hd__xor2_1
XU$$4017 U$$4154/A1 U$$4029/A2 U$$4154/B1 U$$4029/B2 VGND VGND VPWR VPWR U$$4018/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4028 U$$4028/A U$$4044/B VGND VGND VPWR VPWR U$$4028/X sky130_fd_sc_hd__xor2_1
XFILLER_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4039 U$$4176/A1 U$$4071/A2 U$$4176/B1 U$$4071/B2 VGND VGND VPWR VPWR U$$4040/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3305 U$$3305/A U$$3357/B VGND VGND VPWR VPWR U$$3305/X sky130_fd_sc_hd__xor2_1
XU$$3316 U$$3453/A1 U$$3320/A2 U$$3453/B1 U$$3320/B2 VGND VGND VPWR VPWR U$$3317/A
+ sky130_fd_sc_hd__a22o_1
XU$$3327 U$$3327/A U$$3369/B VGND VGND VPWR VPWR U$$3327/X sky130_fd_sc_hd__xor2_1
XU$$3338 U$$4434/A1 U$$3418/A2 U$$4436/A1 U$$3418/B2 VGND VGND VPWR VPWR U$$3339/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3349 U$$3349/A U$$3357/B VGND VGND VPWR VPWR U$$3349/X sky130_fd_sc_hd__xor2_1
XU$$2604 _654_/Q VGND VGND VPWR VPWR U$$2606/B sky130_fd_sc_hd__inv_1
XU$$2615 U$$3024/B1 U$$2663/A2 U$$2754/A1 U$$2663/B2 VGND VGND VPWR VPWR U$$2616/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2626 U$$2626/A U$$2654/B VGND VGND VPWR VPWR U$$2626/X sky130_fd_sc_hd__xor2_1
XFILLER_34_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2637 U$$2909/B1 U$$2687/A2 U$$2774/B1 U$$2687/B2 VGND VGND VPWR VPWR U$$2638/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1903 U$$944/A1 U$$1909/A2 U$$944/B1 U$$1909/B2 VGND VGND VPWR VPWR U$$1904/A sky130_fd_sc_hd__a22o_1
XU$$2648 U$$2648/A U$$2654/B VGND VGND VPWR VPWR U$$2648/X sky130_fd_sc_hd__xor2_1
XU$$2659 U$$330/A1 U$$2663/A2 U$$2796/B1 U$$2663/B2 VGND VGND VPWR VPWR U$$2660/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1914 U$$1914/A U$$1916/B VGND VGND VPWR VPWR U$$1914/X sky130_fd_sc_hd__xor2_1
XU$$1925 U$$1925/A U$$2003/B VGND VGND VPWR VPWR U$$1925/X sky130_fd_sc_hd__xor2_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1936 U$$2895/A1 U$$1976/A2 U$$2210/B1 U$$1976/B2 VGND VGND VPWR VPWR U$$1937/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1947 U$$1947/A U$$2011/B VGND VGND VPWR VPWR U$$1947/X sky130_fd_sc_hd__xor2_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1958 U$$3054/A1 U$$2040/A2 U$$3193/A1 U$$2040/B2 VGND VGND VPWR VPWR U$$1959/A
+ sky130_fd_sc_hd__a22o_1
XU$$1969 U$$1969/A U$$1977/B VGND VGND VPWR VPWR U$$1969/X sky130_fd_sc_hd__xor2_1
XFILLER_148_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1042 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_406_ _559_/CLK _406_/D VGND VGND VPWR VPWR _406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_110 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_337_ _467_/CLK _337_/D VGND VGND VPWR VPWR _337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_268_ _520_/CLK _268_/D VGND VGND VPWR VPWR _268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_199_ _213_/CLK _199_/D VGND VGND VPWR VPWR _199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_71_4 dadda_fa_2_71_4/A dadda_fa_2_71_4/B dadda_fa_2_71_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/CIN dadda_fa_3_71_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_64_3 dadda_fa_2_64_3/A dadda_fa_2_64_3/B dadda_fa_2_64_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/B dadda_fa_3_64_3/B sky130_fd_sc_hd__fa_1
Xrepeater803 U$$2463/B2 VGND VGND VPWR VPWR U$$2423/B2 sky130_fd_sc_hd__buf_4
XFILLER_57_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater814 U$$2197/X VGND VGND VPWR VPWR U$$2318/B2 sky130_fd_sc_hd__buf_4
XFILLER_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater825 U$$2010/B2 VGND VGND VPWR VPWR U$$1982/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_57_2 dadda_fa_2_57_2/A dadda_fa_2_57_2/B dadda_fa_2_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/A dadda_fa_3_57_3/A sky130_fd_sc_hd__fa_1
XFILLER_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater836 U$$1909/B2 VGND VGND VPWR VPWR U$$1915/B2 sky130_fd_sc_hd__buf_6
XFILLER_84_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater847 U$$1553/B2 VGND VGND VPWR VPWR U$$1557/B2 sky130_fd_sc_hd__buf_6
Xrepeater858 U$$263/B2 VGND VGND VPWR VPWR U$$195/B2 sky130_fd_sc_hd__buf_2
Xdadda_fa_5_34_1 dadda_fa_5_34_1/A dadda_fa_5_34_1/B dadda_fa_5_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_35_0/B dadda_fa_7_34_0/A sky130_fd_sc_hd__fa_1
XU$$10 U$$8/B1 U$$8/A2 U$$12/A1 U$$8/B2 VGND VGND VPWR VPWR U$$11/A sky130_fd_sc_hd__a22o_1
Xrepeater869 U$$1478/B2 VGND VGND VPWR VPWR U$$1500/B2 sky130_fd_sc_hd__buf_8
XU$$21 U$$21/A U$$9/B VGND VGND VPWR VPWR U$$21/X sky130_fd_sc_hd__xor2_1
XU$$32 U$$32/A1 U$$68/A2 U$$34/A1 U$$68/B2 VGND VGND VPWR VPWR U$$33/A sky130_fd_sc_hd__a22o_1
XFILLER_37_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$43 U$$43/A U$$57/B VGND VGND VPWR VPWR U$$43/X sky130_fd_sc_hd__xor2_1
XFILLER_64_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_27_0 dadda_fa_5_27_0/A dadda_fa_5_27_0/B dadda_fa_5_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_28_0/A dadda_fa_6_27_0/CIN sky130_fd_sc_hd__fa_1
XU$$54 U$$54/A1 U$$68/A2 U$$56/A1 U$$68/B2 VGND VGND VPWR VPWR U$$55/A sky130_fd_sc_hd__a22o_1
XU$$3850 U$$4259/B1 U$$3874/A2 U$$4400/A1 U$$3874/B2 VGND VGND VPWR VPWR U$$3851/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$65 U$$65/A U$$3/A VGND VGND VPWR VPWR U$$65/X sky130_fd_sc_hd__xor2_1
XU$$76 U$$76/A1 U$$84/A2 U$$78/A1 U$$84/B2 VGND VGND VPWR VPWR U$$77/A sky130_fd_sc_hd__a22o_1
XU$$3861 U$$3861/A U$$3965/B VGND VGND VPWR VPWR U$$3861/X sky130_fd_sc_hd__xor2_1
XU$$87 U$$87/A U$$93/B VGND VGND VPWR VPWR U$$87/X sky130_fd_sc_hd__xor2_1
XU$$3872 _566_/Q U$$3874/A2 U$$584/B1 U$$3874/B2 VGND VGND VPWR VPWR U$$3873/A sky130_fd_sc_hd__a22o_1
XU$$3883 U$$3883/A U$$3917/B VGND VGND VPWR VPWR U$$3883/X sky130_fd_sc_hd__xor2_1
XU$$3894 U$$4442/A1 U$$3910/A2 U$$4031/B1 U$$3910/B2 VGND VGND VPWR VPWR U$$3895/A
+ sky130_fd_sc_hd__a22o_1
XU$$98 U$$98/A1 U$$98/A2 U$$98/B1 U$$98/B2 VGND VGND VPWR VPWR U$$99/A sky130_fd_sc_hd__a22o_1
XFILLER_24_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_12 _278_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_23 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_34 _282_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_45 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_67 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_78 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 _286_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_5_101_0 dadda_fa_5_101_0/A dadda_fa_5_101_0/B dadda_fa_5_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_102_0/A dadda_fa_6_101_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_52_1 U$$776/X U$$909/X U$$1042/X VGND VGND VPWR VPWR dadda_fa_2_53_0/CIN
+ dadda_fa_2_52_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_444 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_45_0 U$$97/X U$$230/X U$$363/X VGND VGND VPWR VPWR dadda_fa_2_46_2/A dadda_fa_2_45_4/B
+ sky130_fd_sc_hd__fa_1
XFILLER_210_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_920 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_56 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_81_3 dadda_fa_3_81_3/A dadda_fa_3_81_3/B dadda_fa_3_81_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_1/B dadda_fa_4_81_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_886 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_74_2 dadda_fa_3_74_2/A dadda_fa_3_74_2/B dadda_fa_3_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_1/A dadda_fa_4_74_2/B sky130_fd_sc_hd__fa_1
XFILLER_3_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_67_1 dadda_fa_3_67_1/A dadda_fa_3_67_1/B dadda_fa_3_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_0/CIN dadda_fa_4_67_2/A sky130_fd_sc_hd__fa_1
XFILLER_78_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_44_0 dadda_fa_6_44_0/A dadda_fa_6_44_0/B dadda_fa_6_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_45_0/B dadda_fa_7_44_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3102 U$$4472/A1 U$$3148/A2 U$$4474/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3103/A
+ sky130_fd_sc_hd__a22o_1
XU$$3113 U$$3113/A U$$3121/B VGND VGND VPWR VPWR U$$3113/X sky130_fd_sc_hd__xor2_1
XU$$3124 U$$3124/A1 U$$3132/A2 U$$3124/B1 U$$3132/B2 VGND VGND VPWR VPWR U$$3125/A
+ sky130_fd_sc_hd__a22o_1
XU$$3135 U$$3135/A U$$3145/B VGND VGND VPWR VPWR U$$3135/X sky130_fd_sc_hd__xor2_1
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2401 U$$3769/B1 U$$2437/A2 U$$3771/B1 U$$2437/B2 VGND VGND VPWR VPWR U$$2402/A
+ sky130_fd_sc_hd__a22o_1
XU$$3146 U$$3283/A1 U$$3018/X U$$3285/A1 U$$3019/X VGND VGND VPWR VPWR U$$3147/A sky130_fd_sc_hd__a22o_1
XFILLER_34_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3157 U$$3157/A1 U$$3209/A2 U$$3157/B1 U$$3209/B2 VGND VGND VPWR VPWR U$$3158/A
+ sky130_fd_sc_hd__a22o_1
XU$$2412 U$$2412/A U$$2436/B VGND VGND VPWR VPWR U$$2412/X sky130_fd_sc_hd__xor2_1
XU$$2423 U$$916/A1 U$$2423/A2 U$$3519/B1 U$$2423/B2 VGND VGND VPWR VPWR U$$2424/A
+ sky130_fd_sc_hd__a22o_1
XU$$3168 U$$3168/A U$$3218/B VGND VGND VPWR VPWR U$$3168/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_103_2 dadda_fa_4_103_2/A dadda_fa_4_103_2/B dadda_fa_4_103_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/CIN dadda_fa_5_103_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2434 U$$2434/A U$$2436/B VGND VGND VPWR VPWR U$$2434/X sky130_fd_sc_hd__xor2_1
XU$$3179 U$$4273/B1 U$$3231/A2 U$$3453/B1 U$$3231/B2 VGND VGND VPWR VPWR U$$3180/A
+ sky130_fd_sc_hd__a22o_1
XU$$1700 U$$467/A1 U$$1718/A2 U$$1976/A1 U$$1718/B2 VGND VGND VPWR VPWR U$$1701/A
+ sky130_fd_sc_hd__a22o_1
XU$$2445 U$$3404/A1 U$$2451/A2 U$$4502/A1 U$$2451/B2 VGND VGND VPWR VPWR U$$2446/A
+ sky130_fd_sc_hd__a22o_1
XU$$1711 U$$1711/A U$$1711/B VGND VGND VPWR VPWR U$$1711/X sky130_fd_sc_hd__xor2_1
XU$$2456 U$$2456/A U$$2462/B VGND VGND VPWR VPWR U$$2456/X sky130_fd_sc_hd__xor2_1
XFILLER_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2467 _652_/Q VGND VGND VPWR VPWR U$$2469/B sky130_fd_sc_hd__inv_1
XU$$1722 U$$761/B1 U$$1740/A2 U$$628/A1 U$$1740/B2 VGND VGND VPWR VPWR U$$1723/A sky130_fd_sc_hd__a22o_1
XU$$1733 U$$1733/A U$$1737/B VGND VGND VPWR VPWR U$$1733/X sky130_fd_sc_hd__xor2_1
XFILLER_15_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2478 U$$2478/A1 U$$2516/A2 U$$3163/B1 U$$2516/B2 VGND VGND VPWR VPWR U$$2479/A
+ sky130_fd_sc_hd__a22o_1
XU$$2489 U$$2489/A U$$2531/B VGND VGND VPWR VPWR U$$2489/X sky130_fd_sc_hd__xor2_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1744 U$$922/A1 U$$1768/A2 U$$924/A1 U$$1768/B2 VGND VGND VPWR VPWR U$$1745/A sky130_fd_sc_hd__a22o_1
XU$$1755 U$$1755/A U$$1763/B VGND VGND VPWR VPWR U$$1755/X sky130_fd_sc_hd__xor2_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1766 U$$944/A1 U$$1768/A2 U$$946/A1 U$$1768/B2 VGND VGND VPWR VPWR U$$1767/A sky130_fd_sc_hd__a22o_1
XFILLER_188_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1777 U$$1777/A U$$1780/A VGND VGND VPWR VPWR U$$1777/X sky130_fd_sc_hd__xor2_1
XFILLER_202_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1788 U$$1788/A U$$1820/B VGND VGND VPWR VPWR U$$1788/X sky130_fd_sc_hd__xor2_1
XU$$1799 U$$18/A1 U$$1851/A2 U$$2210/B1 U$$1851/B2 VGND VGND VPWR VPWR U$$1800/A sky130_fd_sc_hd__a22o_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_117_0 dadda_fa_7_117_0/A dadda_fa_7_117_0/B dadda_fa_7_117_0/CIN VGND
+ VGND VPWR VPWR _542_/D _413_/D sky130_fd_sc_hd__fa_1
XFILLER_174_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput10 a[18] VGND VGND VPWR VPWR _634_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput21 a[28] VGND VGND VPWR VPWR _644_/D sky130_fd_sc_hd__clkbuf_1
Xinput32 a[38] VGND VGND VPWR VPWR _654_/D sky130_fd_sc_hd__clkbuf_1
Xinput43 a[48] VGND VGND VPWR VPWR _664_/D sky130_fd_sc_hd__clkbuf_1
Xinput54 a[58] VGND VGND VPWR VPWR _674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput65 b[0] VGND VGND VPWR VPWR _552_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_200_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput76 b[1] VGND VGND VPWR VPWR _553_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput87 b[2] VGND VGND VPWR VPWR _554_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput98 b[3] VGND VGND VPWR VPWR _555_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater600 U$$1597/A2 VGND VGND VPWR VPWR U$$1553/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_62_0 dadda_fa_2_62_0/A dadda_fa_2_62_0/B dadda_fa_2_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_0/B dadda_fa_3_62_2/B sky130_fd_sc_hd__fa_1
XFILLER_96_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater611 U$$217/A2 VGND VGND VPWR VPWR U$$181/A2 sky130_fd_sc_hd__buf_4
XFILLER_69_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$407 final_adder.U$$324/B final_adder.U$$638/B final_adder.U$$265/X
+ VGND VGND VPWR VPWR final_adder.U$$642/B sky130_fd_sc_hd__a21o_2
XFILLER_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater622 U$$1374/X VGND VGND VPWR VPWR U$$1478/A2 sky130_fd_sc_hd__clkbuf_8
Xfinal_adder.U$$429 final_adder.U$$346/B final_adder.U$$726/B final_adder.U$$309/X
+ VGND VGND VPWR VPWR final_adder.U$$730/B sky130_fd_sc_hd__a21o_2
XFILLER_84_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater633 U$$1176/A2 VGND VGND VPWR VPWR U$$1146/A2 sky130_fd_sc_hd__clkbuf_4
Xrepeater644 U$$964/X VGND VGND VPWR VPWR U$$997/B2 sky130_fd_sc_hd__buf_6
Xrepeater655 U$$827/X VGND VGND VPWR VPWR U$$948/B2 sky130_fd_sc_hd__buf_8
XFILLER_38_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater666 U$$632/B2 VGND VGND VPWR VPWR U$$600/B2 sky130_fd_sc_hd__buf_8
Xrepeater677 U$$4252/X VGND VGND VPWR VPWR U$$4311/B2 sky130_fd_sc_hd__clkbuf_8
Xrepeater688 U$$4115/X VGND VGND VPWR VPWR U$$4226/B2 sky130_fd_sc_hd__buf_4
XFILLER_203_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4370 U$$4370/A U$$4384/A VGND VGND VPWR VPWR U$$4370/X sky130_fd_sc_hd__xor2_1
XFILLER_65_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater699 U$$4065/B2 VGND VGND VPWR VPWR U$$4029/B2 sky130_fd_sc_hd__buf_6
XU$$4381 U$$4516/B1 U$$4381/A2 U$$4381/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4382/A
+ sky130_fd_sc_hd__a22o_1
XU$$4386_1769 VGND VGND VPWR VPWR U$$4386_1769/HI U$$4386/A sky130_fd_sc_hd__conb_1
XFILLER_168_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4392 U$$4392/A1 U$$4388/X U$$4394/A1 U$$4389/X VGND VGND VPWR VPWR U$$4393/A sky130_fd_sc_hd__a22o_1
XFILLER_25_425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3680 U$$3952/B1 U$$3688/A2 U$$4504/A1 U$$3688/B2 VGND VGND VPWR VPWR U$$3681/A
+ sky130_fd_sc_hd__a22o_1
XU$$3691 U$$3691/A U$$3698/A VGND VGND VPWR VPWR U$$3691/X sky130_fd_sc_hd__xor2_1
XFILLER_129_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2990 U$$2990/A U$$3000/B VGND VGND VPWR VPWR U$$2990/X sky130_fd_sc_hd__xor2_1
XFILLER_179_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_439 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_91_2 dadda_fa_4_91_2/A dadda_fa_4_91_2/B dadda_fa_4_91_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_92_0/CIN dadda_fa_5_91_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_193_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_84_1 dadda_fa_4_84_1/A dadda_fa_4_84_1/B dadda_fa_4_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/B dadda_fa_5_84_1/B sky130_fd_sc_hd__fa_1
XFILLER_180_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_61_0 dadda_fa_7_61_0/A dadda_fa_7_61_0/B dadda_fa_7_61_0/CIN VGND VGND
+ VPWR VPWR _486_/D _357_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_77_0 dadda_fa_4_77_0/A dadda_fa_4_77_0/B dadda_fa_4_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/A dadda_fa_5_77_1/A sky130_fd_sc_hd__fa_1
XFILLER_162_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_671_ _679_/CLK _671_/D VGND VGND VPWR VPWR _671_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$802 U$$802/A U$$804/B VGND VGND VPWR VPWR U$$802/X sky130_fd_sc_hd__xor2_1
XFILLER_1_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$813 U$$950/A1 U$$819/A2 U$$950/B1 U$$819/B2 VGND VGND VPWR VPWR U$$814/A sky130_fd_sc_hd__a22o_1
XFILLER_16_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$824 _629_/Q VGND VGND VPWR VPWR U$$824/Y sky130_fd_sc_hd__inv_1
XFILLER_44_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$835 U$$835/A U$$859/B VGND VGND VPWR VPWR U$$835/X sky130_fd_sc_hd__xor2_1
XU$$846 U$$981/B1 U$$878/A2 U$$848/A1 U$$878/B2 VGND VGND VPWR VPWR U$$847/A sky130_fd_sc_hd__a22o_1
XU$$857 U$$857/A U$$935/B VGND VGND VPWR VPWR U$$857/X sky130_fd_sc_hd__xor2_1
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1007 U$$48/A1 U$$979/A2 U$$48/B1 U$$979/B2 VGND VGND VPWR VPWR U$$1008/A sky130_fd_sc_hd__a22o_1
XU$$868 U$$46/A1 U$$878/A2 U$$48/A1 U$$878/B2 VGND VGND VPWR VPWR U$$869/A sky130_fd_sc_hd__a22o_1
XFILLER_16_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$879 U$$879/A U$$879/B VGND VGND VPWR VPWR U$$879/X sky130_fd_sc_hd__xor2_1
XU$$1018 U$$1018/A U$$996/B VGND VGND VPWR VPWR U$$1018/X sky130_fd_sc_hd__xor2_1
XU$$1029 U$$70/A1 U$$999/A2 U$$894/A1 U$$999/B2 VGND VGND VPWR VPWR U$$1030/A sky130_fd_sc_hd__a22o_1
XFILLER_188_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1702 _553_/Q VGND VGND VPWR VPWR U$$4394/A1 sky130_fd_sc_hd__buf_6
XFILLER_137_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_41_5 dadda_fa_2_41_5/A dadda_fa_2_41_5/B dadda_fa_2_41_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_42_2/A dadda_fa_4_41_0/A sky130_fd_sc_hd__fa_2
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_34_4 U$$1937/X U$$2070/X U$$2203/X VGND VGND VPWR VPWR dadda_fa_3_35_1/CIN
+ dadda_fa_3_34_3/CIN sky130_fd_sc_hd__fa_1
XU$$2220 U$$302/A1 U$$2262/A2 U$$989/A1 U$$2262/B2 VGND VGND VPWR VPWR U$$2221/A sky130_fd_sc_hd__a22o_1
XU$$2231 U$$2231/A U$$2243/B VGND VGND VPWR VPWR U$$2231/X sky130_fd_sc_hd__xor2_1
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2242 U$$3884/B1 U$$2242/A2 U$$3751/A1 U$$2242/B2 VGND VGND VPWR VPWR U$$2243/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2253 U$$2253/A U$$2303/B VGND VGND VPWR VPWR U$$2253/X sky130_fd_sc_hd__xor2_1
XFILLER_179_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2264 U$$3769/B1 U$$2274/A2 U$$3771/B1 U$$2274/B2 VGND VGND VPWR VPWR U$$2265/A
+ sky130_fd_sc_hd__a22o_1
XU$$1530 U$$1530/A U$$1558/B VGND VGND VPWR VPWR U$$1530/X sky130_fd_sc_hd__xor2_1
XU$$2275 U$$2275/A U$$2309/B VGND VGND VPWR VPWR U$$2275/X sky130_fd_sc_hd__xor2_1
XU$$1541 U$$2909/B1 U$$1577/A2 U$$2774/B1 U$$1577/B2 VGND VGND VPWR VPWR U$$1542/A
+ sky130_fd_sc_hd__a22o_1
XU$$2286 U$$914/B1 U$$2326/A2 U$$3519/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2287/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2297 U$$2297/A U$$2321/B VGND VGND VPWR VPWR U$$2297/X sky130_fd_sc_hd__xor2_1
XFILLER_22_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1552 U$$1552/A U$$1558/B VGND VGND VPWR VPWR U$$1552/X sky130_fd_sc_hd__xor2_1
XU$$1563 U$$467/A1 U$$1587/A2 U$$3346/A1 U$$1587/B2 VGND VGND VPWR VPWR U$$1564/A
+ sky130_fd_sc_hd__a22o_1
XU$$1574 U$$1574/A U$$1578/B VGND VGND VPWR VPWR U$$1574/X sky130_fd_sc_hd__xor2_1
XFILLER_15_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1585 U$$761/B1 U$$1587/A2 U$$900/B1 U$$1587/B2 VGND VGND VPWR VPWR U$$1586/A sky130_fd_sc_hd__a22o_1
XFILLER_176_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1596 U$$1596/A U$$1598/B VGND VGND VPWR VPWR U$$1596/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_94_0 dadda_fa_5_94_0/A dadda_fa_5_94_0/B dadda_fa_5_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_95_0/A dadda_fa_6_94_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_129_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_79_6 U$$3490/X U$$3623/X U$$3756/X VGND VGND VPWR VPWR dadda_fa_2_80_2/B
+ dadda_fa_2_79_5/B sky130_fd_sc_hd__fa_1
XFILLER_44_1124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$204 final_adder.U$$699/A final_adder.U$$698/A VGND VGND VPWR VPWR
+ final_adder.U$$294/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$215 final_adder.U$$709/A final_adder.U$$581/B1 final_adder.U$$215/B1
+ VGND VGND VPWR VPWR final_adder.U$$215/X sky130_fd_sc_hd__a21o_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$226 final_adder.U$$721/A final_adder.U$$720/A VGND VGND VPWR VPWR
+ final_adder.U$$304/A sky130_fd_sc_hd__and2_1
Xrepeater430 U$$415/X VGND VGND VPWR VPWR U$$545/A2 sky130_fd_sc_hd__clkbuf_8
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater441 U$$62/A2 VGND VGND VPWR VPWR U$$68/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$237 final_adder.U$$731/A final_adder.U$$603/B1 final_adder.U$$237/B1
+ VGND VGND VPWR VPWR final_adder.U$$237/X sky130_fd_sc_hd__a21o_1
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$248 final_adder.U$$743/A final_adder.U$$742/A VGND VGND VPWR VPWR
+ final_adder.U$$316/B sky130_fd_sc_hd__and2_1
Xrepeater452 U$$3977/X VGND VGND VPWR VPWR U$$4095/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$259 final_adder.U$$258/A final_adder.U$$133/X final_adder.U$$135/X
+ VGND VGND VPWR VPWR final_adder.U$$259/X sky130_fd_sc_hd__a21o_1
Xrepeater463 U$$3823/A2 VGND VGND VPWR VPWR U$$3769/A2 sky130_fd_sc_hd__buf_6
XU$$109 U$$109/A U$$117/B VGND VGND VPWR VPWR U$$109/X sky130_fd_sc_hd__xor2_1
XFILLER_26_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater474 U$$3674/A2 VGND VGND VPWR VPWR U$$3688/A2 sky130_fd_sc_hd__buf_6
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater485 U$$3429/X VGND VGND VPWR VPWR U$$3555/A2 sky130_fd_sc_hd__buf_6
Xrepeater496 U$$3231/A2 VGND VGND VPWR VPWR U$$3215/A2 sky130_fd_sc_hd__buf_4
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$682_1842 VGND VGND VPWR VPWR U$$682_1842/HI U$$682/B1 sky130_fd_sc_hd__conb_1
XFILLER_26_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1009 U$$2843/B VGND VGND VPWR VPWR U$$2875/B sky130_fd_sc_hd__buf_6
XFILLER_181_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_110_2 U$$3951/X U$$4084/X U$$4217/X VGND VGND VPWR VPWR dadda_fa_4_111_1/B
+ dadda_fa_4_110_2/B sky130_fd_sc_hd__fa_1
XFILLER_119_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_103_1 U$$4336/X U$$4469/X input133/X VGND VGND VPWR VPWR dadda_fa_4_104_0/CIN
+ dadda_fa_4_103_2/A sky130_fd_sc_hd__fa_1
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_558 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput200 c[49] VGND VGND VPWR VPWR input200/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput211 c[59] VGND VGND VPWR VPWR input211/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_124_0 dadda_fa_6_124_0/A dadda_fa_6_124_0/B dadda_fa_6_124_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_125_0/B dadda_fa_7_124_0/CIN sky130_fd_sc_hd__fa_1
Xinput222 c[69] VGND VGND VPWR VPWR input222/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput233 c[79] VGND VGND VPWR VPWR input233/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput244 c[89] VGND VGND VPWR VPWR input244/X sky130_fd_sc_hd__buf_2
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_494 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_67_4 U$$1737/X U$$1870/X U$$2003/X VGND VGND VPWR VPWR dadda_fa_1_68_6/CIN
+ dadda_fa_1_67_8/CIN sky130_fd_sc_hd__fa_1
Xdadda_ha_3_116_0_1876 VGND VGND VPWR VPWR dadda_ha_3_116_0/A dadda_ha_3_116_0_1876/LO
+ sky130_fd_sc_hd__conb_1
Xinput255 c[99] VGND VGND VPWR VPWR input255/X sky130_fd_sc_hd__buf_4
XTAP_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_44_3 dadda_fa_3_44_3/A dadda_fa_3_44_3/B dadda_fa_3_44_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_1/B dadda_fa_4_44_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$610 U$$882/B1 U$$616/A2 U$$747/B1 U$$616/B2 VGND VGND VPWR VPWR U$$611/A sky130_fd_sc_hd__a22o_1
X_654_ _662_/CLK _654_/D VGND VGND VPWR VPWR _654_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_37_2 dadda_fa_3_37_2/A dadda_fa_3_37_2/B dadda_fa_3_37_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_1/A dadda_fa_4_37_2/B sky130_fd_sc_hd__fa_1
XU$$621 U$$621/A U$$665/B VGND VGND VPWR VPWR U$$621/X sky130_fd_sc_hd__xor2_1
XU$$632 U$$84/A1 U$$632/A2 U$$84/B1 U$$632/B2 VGND VGND VPWR VPWR U$$633/A sky130_fd_sc_hd__a22o_1
XU$$643 U$$643/A U$$651/B VGND VGND VPWR VPWR U$$643/X sky130_fd_sc_hd__xor2_1
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$654 U$$791/A1 U$$682/A2 U$$791/B1 U$$682/B2 VGND VGND VPWR VPWR U$$655/A sky130_fd_sc_hd__a22o_1
XFILLER_1_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1003 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_585_ _588_/CLK _585_/D VGND VGND VPWR VPWR _585_/Q sky130_fd_sc_hd__dfxtp_1
XU$$665 U$$665/A U$$665/B VGND VGND VPWR VPWR U$$665/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$676 U$$676/A1 U$$682/A2 U$$676/B1 U$$682/B2 VGND VGND VPWR VPWR U$$677/A sky130_fd_sc_hd__a22o_1
XFILLER_186_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$687 U$$810/B VGND VGND VPWR VPWR U$$687/Y sky130_fd_sc_hd__inv_1
XFILLER_140_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$698 U$$698/A U$$726/B VGND VGND VPWR VPWR U$$698/X sky130_fd_sc_hd__xor2_1
XFILLER_108_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1510 U$$56/A1 VGND VGND VPWR VPWR U$$330/A1 sky130_fd_sc_hd__buf_4
XFILLER_67_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1521 U$$3342/A1 VGND VGND VPWR VPWR U$$54/A1 sky130_fd_sc_hd__buf_4
XFILLER_193_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1532 _573_/Q VGND VGND VPWR VPWR U$$4434/A1 sky130_fd_sc_hd__buf_4
Xrepeater1543 U$$2786/B1 VGND VGND VPWR VPWR U$$596/A1 sky130_fd_sc_hd__buf_4
XFILLER_158_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1554 U$$4154/B1 VGND VGND VPWR VPWR U$$4293/A1 sky130_fd_sc_hd__buf_6
Xrepeater1565 U$$3193/A1 VGND VGND VPWR VPWR U$$42/A1 sky130_fd_sc_hd__buf_6
XFILLER_181_992 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_89_5 dadda_fa_2_89_5/A dadda_fa_2_89_5/B dadda_fa_2_89_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_90_2/A dadda_fa_4_89_0/A sky130_fd_sc_hd__fa_2
XFILLER_119_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1576 U$$4287/A1 VGND VGND VPWR VPWR U$$2641/B1 sky130_fd_sc_hd__buf_4
XFILLER_4_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1587 U$$310/A1 VGND VGND VPWR VPWR U$$582/B1 sky130_fd_sc_hd__buf_6
XFILLER_165_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1598 U$$4007/A1 VGND VGND VPWR VPWR U$$3320/B1 sky130_fd_sc_hd__buf_4
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4417_1787 VGND VGND VPWR VPWR U$$4417_1787/HI U$$4417/B sky130_fd_sc_hd__conb_1
XFILLER_119_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_26_2 U$$857/X U$$990/X VGND VGND VPWR VPWR dadda_fa_3_27_3/A dadda_fa_4_26_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_95_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_32_1 U$$470/X U$$603/X U$$736/X VGND VGND VPWR VPWR dadda_fa_3_33_0/CIN
+ dadda_fa_3_32_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_1204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2050 U$$2459/B1 U$$2052/A2 U$$2872/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2051/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_25_0 U$$57/X U$$190/X U$$323/X VGND VGND VPWR VPWR dadda_fa_3_26_2/CIN
+ dadda_fa_3_25_3/CIN sky130_fd_sc_hd__fa_1
XU$$2061 U$$2061/A1 U$$2129/A2 U$$2746/B1 U$$2129/B2 VGND VGND VPWR VPWR U$$2062/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2072 U$$2072/A U$$2108/B VGND VGND VPWR VPWR U$$2072/X sky130_fd_sc_hd__xor2_1
XFILLER_35_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2083 U$$302/A1 U$$2129/A2 U$$989/A1 U$$2129/B2 VGND VGND VPWR VPWR U$$2084/A sky130_fd_sc_hd__a22o_1
XU$$2094 U$$2094/A U$$2144/B VGND VGND VPWR VPWR U$$2094/X sky130_fd_sc_hd__xor2_1
XFILLER_200_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1360 U$$1360/A U$$1368/B VGND VGND VPWR VPWR U$$1360/X sky130_fd_sc_hd__xor2_1
XU$$1371 _636_/Q VGND VGND VPWR VPWR U$$1373/B sky130_fd_sc_hd__inv_1
XU$$1382 U$$2613/B1 U$$1424/A2 U$$562/A1 U$$1424/B2 VGND VGND VPWR VPWR U$$1383/A
+ sky130_fd_sc_hd__a22o_1
XU$$1393 U$$1393/A U$$1459/B VGND VGND VPWR VPWR U$$1393/X sky130_fd_sc_hd__xor2_1
XFILLER_200_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_119_1 dadda_fa_5_119_1/A dadda_fa_5_119_1/B dadda_fa_5_119_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_120_0/B dadda_fa_7_119_0/A sky130_fd_sc_hd__fa_1
XFILLER_191_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_84_4 U$$2968/X U$$3101/X U$$3234/X VGND VGND VPWR VPWR dadda_fa_2_85_3/B
+ dadda_fa_2_84_5/B sky130_fd_sc_hd__fa_1
XFILLER_116_396 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_77_3 U$$2555/X U$$2688/X U$$2821/X VGND VGND VPWR VPWR dadda_fa_2_78_1/B
+ dadda_fa_2_77_4/B sky130_fd_sc_hd__fa_1
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_54_2 dadda_fa_4_54_2/A dadda_fa_4_54_2/B dadda_fa_4_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/CIN dadda_fa_5_54_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_47_1 dadda_fa_4_47_1/A dadda_fa_4_47_1/B dadda_fa_4_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/B dadda_fa_5_47_1/B sky130_fd_sc_hd__fa_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_24_0 dadda_fa_7_24_0/A dadda_fa_7_24_0/B dadda_fa_7_24_0/CIN VGND VGND
+ VPWR VPWR _449_/D _320_/D sky130_fd_sc_hd__fa_1
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_305 _235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_316 _237_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_327 _239_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 U$$785/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_349 U$$896/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_370_ _500_/CLK _370_/D VGND VGND VPWR VPWR _370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_926 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_72_2 U$$1348/X U$$1481/X U$$1614/X VGND VGND VPWR VPWR dadda_fa_1_73_7/CIN
+ dadda_fa_1_72_8/CIN sky130_fd_sc_hd__fa_1
XTAP_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_65_1 U$$536/X U$$669/X U$$802/X VGND VGND VPWR VPWR dadda_fa_1_66_5/CIN
+ dadda_fa_1_65_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_77_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_42_0 dadda_fa_3_42_0/A dadda_fa_3_42_0/B dadda_fa_3_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_0/B dadda_fa_4_42_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_58_0 U$$123/X U$$256/X U$$389/X VGND VGND VPWR VPWR dadda_fa_1_59_6/CIN
+ dadda_fa_1_58_8/A sky130_fd_sc_hd__fa_1
XTAP_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$440 U$$440/A U$$456/B VGND VGND VPWR VPWR U$$440/X sky130_fd_sc_hd__xor2_1
X_637_ _637_/CLK _637_/D VGND VGND VPWR VPWR _637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_478 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$451 U$$451/A1 U$$499/A2 U$$999/B1 U$$499/B2 VGND VGND VPWR VPWR U$$452/A sky130_fd_sc_hd__a22o_1
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$462 U$$462/A U$$532/B VGND VGND VPWR VPWR U$$462/X sky130_fd_sc_hd__xor2_1
XU$$473 U$$882/B1 U$$483/A2 U$$747/B1 U$$483/B2 VGND VGND VPWR VPWR U$$474/A sky130_fd_sc_hd__a22o_1
XFILLER_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$484 U$$484/A U$$484/B VGND VGND VPWR VPWR U$$484/X sky130_fd_sc_hd__xor2_1
XFILLER_204_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_568_ _569_/CLK _568_/D VGND VGND VPWR VPWR _568_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$495 U$$84/A1 U$$499/A2 U$$84/B1 U$$499/B2 VGND VGND VPWR VPWR U$$496/A sky130_fd_sc_hd__a22o_1
XFILLER_44_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_499_ _500_/CLK _499_/D VGND VGND VPWR VPWR _499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_94_3 U$$3919/X U$$4052/X U$$4185/X VGND VGND VPWR VPWR dadda_fa_3_95_1/B
+ dadda_fa_3_94_3/B sky130_fd_sc_hd__fa_1
XFILLER_145_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1340 U$$3521/B1 VGND VGND VPWR VPWR U$$781/B1 sky130_fd_sc_hd__buf_4
XFILLER_154_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1351 U$$3658/A1 VGND VGND VPWR VPWR U$$3932/A1 sky130_fd_sc_hd__buf_6
XFILLER_172_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1362 _595_/Q VGND VGND VPWR VPWR U$$3791/B1 sky130_fd_sc_hd__buf_6
XFILLER_126_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_87_2 U$$4437/X input242/X dadda_fa_2_87_2/CIN VGND VGND VPWR VPWR dadda_fa_3_88_1/A
+ dadda_fa_3_87_3/A sky130_fd_sc_hd__fa_1
Xrepeater1373 U$$3652/A1 VGND VGND VPWR VPWR U$$912/A1 sky130_fd_sc_hd__buf_4
Xrepeater1384 _592_/Q VGND VGND VPWR VPWR U$$4061/A1 sky130_fd_sc_hd__buf_4
XFILLER_114_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_64_1 dadda_fa_5_64_1/A dadda_fa_5_64_1/B dadda_fa_5_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_65_0/B dadda_fa_7_64_0/A sky130_fd_sc_hd__fa_1
XFILLER_99_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1395 U$$3783/A1 VGND VGND VPWR VPWR U$$906/A1 sky130_fd_sc_hd__buf_4
XFILLER_141_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_57_0 dadda_fa_5_57_0/A dadda_fa_5_57_0/B dadda_fa_5_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_58_0/A dadda_fa_6_57_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_56_8 dadda_fa_1_56_8/A dadda_fa_1_56_8/B dadda_fa_1_56_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_57_3/A dadda_fa_3_56_0/A sky130_fd_sc_hd__fa_2
XFILLER_41_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_103_0 U$$2739/Y U$$2873/X U$$3006/X VGND VGND VPWR VPWR dadda_fa_3_104_2/B
+ dadda_fa_3_103_3/B sky130_fd_sc_hd__fa_1
XFILLER_39_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1190 U$$94/A1 U$$1190/A2 U$$96/A1 U$$1190/B2 VGND VGND VPWR VPWR U$$1191/A sky130_fd_sc_hd__a22o_1
XFILLER_206_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_723 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1043 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_82_1 U$$1634/X U$$1767/X U$$1900/X VGND VGND VPWR VPWR dadda_fa_2_83_1/CIN
+ dadda_fa_2_82_4/A sky130_fd_sc_hd__fa_1
XFILLER_172_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_75_0 U$$1620/X U$$1753/X U$$1886/X VGND VGND VPWR VPWR dadda_fa_2_76_0/B
+ dadda_fa_2_75_3/B sky130_fd_sc_hd__fa_1
XFILLER_137_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3509 U$$3646/A1 U$$3429/X U$$4470/A1 U$$3430/X VGND VGND VPWR VPWR U$$3510/A sky130_fd_sc_hd__a22o_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2808 U$$4176/B1 U$$2832/A2 U$$3495/A1 U$$2832/B2 VGND VGND VPWR VPWR U$$2809/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2819 U$$2819/A U$$2861/B VGND VGND VPWR VPWR U$$2819/X sky130_fd_sc_hd__xor2_1
XANTENNA_102 _287_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _290_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_146 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _180_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_422_ _627_/CLK _422_/D VGND VGND VPWR VPWR _422_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _183_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_179 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_353_ _353_/CLK _353_/D VGND VGND VPWR VPWR _353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_284_ _526_/CLK _284_/D VGND VGND VPWR VPWR _284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_97_1 dadda_fa_3_97_1/A dadda_fa_3_97_1/B dadda_fa_3_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_0/CIN dadda_fa_4_97_2/A sky130_fd_sc_hd__fa_1
XFILLER_5_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_74_0 dadda_fa_6_74_0/A dadda_fa_6_74_0/B dadda_fa_6_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_75_0/B dadda_fa_7_74_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1043 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 a[16] VGND VGND VPWR VPWR _632_/D sky130_fd_sc_hd__clkbuf_2
XTAP_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_119_0 U$$3835/Y U$$3969/X U$$4102/X VGND VGND VPWR VPWR dadda_fa_5_120_0/CIN
+ dadda_fa_5_119_1/B sky130_fd_sc_hd__fa_1
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$270 U$$270/A U$$272/B VGND VGND VPWR VPWR U$$270/X sky130_fd_sc_hd__xor2_1
XFILLER_33_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$281 U$$281/A U$$319/B VGND VGND VPWR VPWR U$$281/X sky130_fd_sc_hd__xor2_1
XU$$292 U$$429/A1 U$$308/A2 U$$429/B1 U$$308/B2 VGND VGND VPWR VPWR U$$293/A sky130_fd_sc_hd__a22o_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$6 _430_/Q _302_/Q VGND VGND VPWR VPWR final_adder.U$$6/COUT final_adder.U$$628/A
+ sky130_fd_sc_hd__ha_1
XFILLER_134_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1038 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput301 _192_/Q VGND VGND VPWR VPWR o[24] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_0 U$$2984/X U$$3117/X U$$3250/X VGND VGND VPWR VPWR dadda_fa_3_93_0/B
+ dadda_fa_3_92_2/B sky130_fd_sc_hd__fa_1
XFILLER_145_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput312 _202_/Q VGND VGND VPWR VPWR o[34] sky130_fd_sc_hd__buf_2
XFILLER_195_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput323 _212_/Q VGND VGND VPWR VPWR o[44] sky130_fd_sc_hd__buf_2
XFILLER_173_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput334 _222_/Q VGND VGND VPWR VPWR o[54] sky130_fd_sc_hd__buf_2
Xoutput345 _232_/Q VGND VGND VPWR VPWR o[64] sky130_fd_sc_hd__buf_2
Xoutput356 _242_/Q VGND VGND VPWR VPWR o[74] sky130_fd_sc_hd__buf_2
Xrepeater1170 U$$410/A VGND VGND VPWR VPWR U$$393/B sky130_fd_sc_hd__buf_6
Xoutput367 _252_/Q VGND VGND VPWR VPWR o[84] sky130_fd_sc_hd__buf_2
Xrepeater1181 _619_/Q VGND VGND VPWR VPWR U$$272/B sky130_fd_sc_hd__buf_4
XFILLER_114_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput378 _262_/Q VGND VGND VPWR VPWR o[94] sky130_fd_sc_hd__buf_2
XFILLER_160_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1192 U$$4105/B1 VGND VGND VPWR VPWR U$$406/B1 sky130_fd_sc_hd__buf_4
Xdadda_ha_4_118_2 U$$4499/X input149/X VGND VGND VPWR VPWR dadda_fa_5_119_1/A dadda_ha_4_118_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_141_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_6 dadda_fa_1_61_6/A dadda_fa_1_61_6/B dadda_fa_1_61_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_2/B dadda_fa_2_61_5/B sky130_fd_sc_hd__fa_1
XFILLER_45_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_54_5 U$$2775/X U$$2908/X U$$3041/X VGND VGND VPWR VPWR dadda_fa_2_55_2/A
+ dadda_fa_2_54_5/A sky130_fd_sc_hd__fa_1
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_47_4 U$$1697/X U$$1830/X U$$1963/X VGND VGND VPWR VPWR dadda_fa_2_48_2/CIN
+ dadda_fa_2_47_5/B sky130_fd_sc_hd__fa_1
XFILLER_55_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_17_2 dadda_fa_4_17_2/A dadda_fa_4_17_2/B dadda_ha_3_17_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_18_0/CIN dadda_fa_5_17_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_91_0 dadda_fa_7_91_0/A dadda_fa_7_91_0/B dadda_fa_7_91_0/CIN VGND VGND
+ VPWR VPWR _516_/D _387_/D sky130_fd_sc_hd__fa_2
XFILLER_137_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4007 U$$4007/A1 U$$4065/A2 _566_/Q U$$4065/B2 VGND VGND VPWR VPWR U$$4008/A sky130_fd_sc_hd__a22o_1
XU$$4018 U$$4018/A U$$4058/B VGND VGND VPWR VPWR U$$4018/X sky130_fd_sc_hd__xor2_1
XFILLER_120_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4029 U$$4440/A1 U$$4029/A2 U$$4442/A1 U$$4029/B2 VGND VGND VPWR VPWR U$$4030/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3306 U$$3578/B1 U$$3356/A2 U$$3445/A1 U$$3356/B2 VGND VGND VPWR VPWR U$$3307/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3317 U$$3317/A U$$3343/B VGND VGND VPWR VPWR U$$3317/X sky130_fd_sc_hd__xor2_1
XU$$3328 U$$3602/A1 U$$3368/A2 U$$4426/A1 U$$3368/B2 VGND VGND VPWR VPWR U$$3329/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3339 U$$3339/A U$$3424/A VGND VGND VPWR VPWR U$$3339/X sky130_fd_sc_hd__xor2_1
XFILLER_73_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2605 _655_/Q VGND VGND VPWR VPWR U$$2605/Y sky130_fd_sc_hd__inv_1
XU$$2616 U$$2616/A U$$2664/B VGND VGND VPWR VPWR U$$2616/X sky130_fd_sc_hd__xor2_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2627 U$$3584/B1 U$$2653/A2 U$$3451/A1 U$$2653/B2 VGND VGND VPWR VPWR U$$2628/A
+ sky130_fd_sc_hd__a22o_1
XU$$2638 U$$2638/A U$$2688/B VGND VGND VPWR VPWR U$$2638/X sky130_fd_sc_hd__xor2_1
XFILLER_46_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1904 U$$1904/A U$$1916/B VGND VGND VPWR VPWR U$$1904/X sky130_fd_sc_hd__xor2_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2649 U$$866/B1 U$$2653/A2 U$$2786/B1 U$$2653/B2 VGND VGND VPWR VPWR U$$2650/A
+ sky130_fd_sc_hd__a22o_1
XU$$1915 U$$817/B1 U$$1915/A2 U$$1915/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1916/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1926 U$$967/A1 U$$1922/X U$$969/A1 U$$1923/X VGND VGND VPWR VPWR U$$1927/A sky130_fd_sc_hd__a22o_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1937 U$$1937/A U$$1977/B VGND VGND VPWR VPWR U$$1937/X sky130_fd_sc_hd__xor2_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1948 U$$2494/B1 U$$1956/A2 U$$854/A1 U$$1956/B2 VGND VGND VPWR VPWR U$$1949/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1959 U$$1959/A U$$2043/B VGND VGND VPWR VPWR U$$1959/X sky130_fd_sc_hd__xor2_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_405_ _534_/CLK _405_/D VGND VGND VPWR VPWR _405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_336_ _466_/CLK _336_/D VGND VGND VPWR VPWR _336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_267_ _520_/CLK _267_/D VGND VGND VPWR VPWR _267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_198_ _213_/CLK _198_/D VGND VGND VPWR VPWR _198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_71_5 dadda_fa_2_71_5/A dadda_fa_2_71_5/B dadda_fa_2_71_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_2/A dadda_fa_4_71_0/A sky130_fd_sc_hd__fa_1
XFILLER_111_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_280 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_64_4 dadda_fa_2_64_4/A dadda_fa_2_64_4/B dadda_fa_2_64_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/CIN dadda_fa_3_64_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater804 U$$2451/B2 VGND VGND VPWR VPWR U$$2463/B2 sky130_fd_sc_hd__buf_6
Xrepeater815 U$$2135/B2 VGND VGND VPWR VPWR U$$2129/B2 sky130_fd_sc_hd__buf_4
Xrepeater826 U$$2038/B2 VGND VGND VPWR VPWR U$$2010/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_57_3 dadda_fa_2_57_3/A dadda_fa_2_57_3/B dadda_fa_2_57_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/B dadda_fa_3_57_3/B sky130_fd_sc_hd__fa_1
Xrepeater837 U$$1907/B2 VGND VGND VPWR VPWR U$$1909/B2 sky130_fd_sc_hd__buf_6
XFILLER_111_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater848 U$$1597/B2 VGND VGND VPWR VPWR U$$1553/B2 sky130_fd_sc_hd__buf_4
XFILLER_49_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$11 U$$11/A U$$9/B VGND VGND VPWR VPWR U$$11/X sky130_fd_sc_hd__xor2_1
Xrepeater859 U$$217/B2 VGND VGND VPWR VPWR U$$181/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$22 U$$22/A1 U$$52/A2 U$$22/B1 U$$52/B2 VGND VGND VPWR VPWR U$$23/A sky130_fd_sc_hd__a22o_1
XU$$33 U$$33/A U$$57/B VGND VGND VPWR VPWR U$$33/X sky130_fd_sc_hd__xor2_1
XFILLER_92_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$44 U$$44/A1 U$$52/A2 U$$46/A1 U$$52/B2 VGND VGND VPWR VPWR U$$45/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_27_1 dadda_fa_5_27_1/A dadda_fa_5_27_1/B dadda_fa_5_27_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_28_0/B dadda_fa_7_27_0/A sky130_fd_sc_hd__fa_2
XU$$55 U$$55/A U$$57/B VGND VGND VPWR VPWR U$$55/X sky130_fd_sc_hd__xor2_1
XU$$3840 U$$3838/Y _672_/Q U$$3836/A U$$3839/X U$$3836/Y VGND VGND VPWR VPWR U$$3840/X
+ sky130_fd_sc_hd__a32o_4
XU$$66 U$$66/A1 U$$68/A2 U$$66/B1 U$$68/B2 VGND VGND VPWR VPWR U$$67/A sky130_fd_sc_hd__a22o_1
XFILLER_64_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3851 U$$3851/A U$$3873/B VGND VGND VPWR VPWR U$$3851/X sky130_fd_sc_hd__xor2_1
XFILLER_25_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3862 U$$4273/A1 U$$3970/A2 U$$4136/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3863/A
+ sky130_fd_sc_hd__a22o_1
XU$$77 U$$77/A U$$81/B VGND VGND VPWR VPWR U$$77/X sky130_fd_sc_hd__xor2_1
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3873 U$$3873/A U$$3873/B VGND VGND VPWR VPWR U$$3873/X sky130_fd_sc_hd__xor2_1
XU$$88 U$$88/A1 U$$4/X U$$90/A1 U$$5/X VGND VGND VPWR VPWR U$$89/A sky130_fd_sc_hd__a22o_1
XFILLER_80_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3884 U$$4156/B1 U$$3916/A2 U$$3884/B1 U$$3916/B2 VGND VGND VPWR VPWR U$$3885/A
+ sky130_fd_sc_hd__a22o_1
XU$$99 U$$99/A U$$99/B VGND VGND VPWR VPWR U$$99/X sky130_fd_sc_hd__xor2_1
XFILLER_197_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_448 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3895 U$$3895/A U$$3895/B VGND VGND VPWR VPWR U$$3895/X sky130_fd_sc_hd__xor2_1
XFILLER_178_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_13 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_24 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_35 _282_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_79 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1097 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_101_1 dadda_fa_5_101_1/A dadda_fa_5_101_1/B dadda_fa_5_101_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_102_0/B dadda_fa_7_101_0/A sky130_fd_sc_hd__fa_2
XFILLER_173_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_39_2 U$$883/X U$$1016/X VGND VGND VPWR VPWR dadda_fa_2_40_4/CIN dadda_fa_3_39_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_56_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_52_2 U$$1175/X U$$1308/X U$$1441/X VGND VGND VPWR VPWR dadda_fa_2_53_1/A
+ dadda_fa_2_52_4/A sky130_fd_sc_hd__fa_1
XFILLER_29_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_45_1 U$$496/X U$$629/X U$$762/X VGND VGND VPWR VPWR dadda_fa_2_46_2/B
+ dadda_fa_2_45_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_22_0 dadda_fa_4_22_0/A dadda_fa_4_22_0/B dadda_fa_4_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/A dadda_fa_5_22_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_38_0 U$$83/X U$$216/X U$$349/X VGND VGND VPWR VPWR dadda_fa_2_39_4/B dadda_fa_2_38_5/B
+ sky130_fd_sc_hd__fa_1
XFILLER_15_139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_278 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_976 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_898 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_74_3 dadda_fa_3_74_3/A dadda_fa_3_74_3/B dadda_fa_3_74_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_1/B dadda_fa_4_74_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_67_2 dadda_fa_3_67_2/A dadda_fa_3_67_2/B dadda_fa_3_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_1/A dadda_fa_4_67_2/B sky130_fd_sc_hd__fa_1
XFILLER_152_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_37_0 dadda_fa_6_37_0/A dadda_fa_6_37_0/B dadda_fa_6_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_38_0/B dadda_fa_7_37_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3103 U$$3103/A U$$3107/B VGND VGND VPWR VPWR U$$3103/X sky130_fd_sc_hd__xor2_1
XFILLER_207_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3114 U$$3934/B1 U$$3132/A2 U$$3799/B1 U$$3132/B2 VGND VGND VPWR VPWR U$$3115/A
+ sky130_fd_sc_hd__a22o_1
XU$$3125 U$$3125/A U$$3133/B VGND VGND VPWR VPWR U$$3125/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3136 U$$3273/A1 U$$3144/A2 U$$3412/A1 U$$3144/B2 VGND VGND VPWR VPWR U$$3137/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2402 U$$2402/A U$$2442/B VGND VGND VPWR VPWR U$$2402/X sky130_fd_sc_hd__xor2_1
XFILLER_46_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3147 U$$3147/A _661_/Q VGND VGND VPWR VPWR U$$3147/X sky130_fd_sc_hd__xor2_1
XU$$2413 U$$3096/B1 U$$2435/A2 U$$2415/A1 U$$2435/B2 VGND VGND VPWR VPWR U$$2414/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3158 U$$3158/A U$$3208/B VGND VGND VPWR VPWR U$$3158/X sky130_fd_sc_hd__xor2_1
XU$$2424 U$$2424/A U$$2462/B VGND VGND VPWR VPWR U$$2424/X sky130_fd_sc_hd__xor2_1
XU$$3169 U$$3578/B1 U$$3215/A2 U$$3445/A1 U$$3215/B2 VGND VGND VPWR VPWR U$$3170/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2435 U$$2435/A1 U$$2435/A2 U$$791/B1 U$$2435/B2 VGND VGND VPWR VPWR U$$2436/A
+ sky130_fd_sc_hd__a22o_1
XU$$1701 U$$1701/A U$$1719/B VGND VGND VPWR VPWR U$$1701/X sky130_fd_sc_hd__xor2_1
XU$$2446 U$$2446/A U$$2466/A VGND VGND VPWR VPWR U$$2446/X sky130_fd_sc_hd__xor2_1
XU$$1712 U$$3354/B1 U$$1762/A2 U$$3221/A1 U$$1762/B2 VGND VGND VPWR VPWR U$$1713/A
+ sky130_fd_sc_hd__a22o_1
XU$$2457 _612_/Q U$$2463/A2 U$$2459/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2458/A sky130_fd_sc_hd__a22o_1
XFILLER_62_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2468 _653_/Q VGND VGND VPWR VPWR U$$2468/Y sky130_fd_sc_hd__inv_1
XU$$1723 U$$1723/A U$$1723/B VGND VGND VPWR VPWR U$$1723/X sky130_fd_sc_hd__xor2_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1734 U$$4474/A1 U$$1648/X U$$92/A1 U$$1649/X VGND VGND VPWR VPWR U$$1735/A sky130_fd_sc_hd__a22o_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2479 U$$2479/A U$$2541/B VGND VGND VPWR VPWR U$$2479/X sky130_fd_sc_hd__xor2_1
XU$$1745 U$$1745/A U$$1747/B VGND VGND VPWR VPWR U$$1745/X sky130_fd_sc_hd__xor2_1
XU$$1756 U$$3124/B1 U$$1762/A2 U$$2991/A1 U$$1762/B2 VGND VGND VPWR VPWR U$$1757/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1767 U$$1767/A U$$1773/B VGND VGND VPWR VPWR U$$1767/X sky130_fd_sc_hd__xor2_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1778 U$$545/A1 U$$1778/A2 U$$1778/B1 U$$1778/B2 VGND VGND VPWR VPWR U$$1779/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1789 U$$967/A1 U$$1859/A2 U$$969/A1 U$$1859/B2 VGND VGND VPWR VPWR U$$1790/A sky130_fd_sc_hd__a22o_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_319_ _448_/CLK _319_/D VGND VGND VPWR VPWR _319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput11 a[19] VGND VGND VPWR VPWR _635_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 a[29] VGND VGND VPWR VPWR _645_/D sky130_fd_sc_hd__clkbuf_1
Xinput33 a[39] VGND VGND VPWR VPWR _655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput44 a[49] VGND VGND VPWR VPWR _665_/D sky130_fd_sc_hd__clkbuf_1
Xinput55 a[59] VGND VGND VPWR VPWR _675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput66 b[10] VGND VGND VPWR VPWR _562_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput77 b[20] VGND VGND VPWR VPWR _572_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput88 b[30] VGND VGND VPWR VPWR _582_/D sky130_fd_sc_hd__clkbuf_1
Xinput99 b[40] VGND VGND VPWR VPWR _592_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_62_1 dadda_fa_2_62_1/A dadda_fa_2_62_1/B dadda_fa_2_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_0/CIN dadda_fa_3_62_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater601 U$$1607/A2 VGND VGND VPWR VPWR U$$1597/A2 sky130_fd_sc_hd__buf_4
XFILLER_96_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater612 U$$217/A2 VGND VGND VPWR VPWR U$$249/A2 sky130_fd_sc_hd__buf_6
XFILLER_57_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$419 final_adder.U$$336/B final_adder.U$$686/B final_adder.U$$289/X
+ VGND VGND VPWR VPWR final_adder.U$$690/B sky130_fd_sc_hd__a21o_2
Xrepeater623 U$$1374/X VGND VGND VPWR VPWR U$$1474/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_55_0 dadda_fa_2_55_0/A dadda_fa_2_55_0/B dadda_fa_2_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_0/B dadda_fa_3_55_2/B sky130_fd_sc_hd__fa_1
Xrepeater634 U$$1190/A2 VGND VGND VPWR VPWR U$$1176/A2 sky130_fd_sc_hd__buf_4
Xrepeater645 U$$1093/B2 VGND VGND VPWR VPWR U$$1089/B2 sky130_fd_sc_hd__buf_4
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater656 U$$765/B2 VGND VGND VPWR VPWR U$$747/B2 sky130_fd_sc_hd__buf_4
Xrepeater667 U$$622/B2 VGND VGND VPWR VPWR U$$632/B2 sky130_fd_sc_hd__buf_8
XU$$4360 U$$4360/A U$$4382/B VGND VGND VPWR VPWR U$$4360/X sky130_fd_sc_hd__xor2_1
Xrepeater678 U$$4252/X VGND VGND VPWR VPWR U$$4345/B2 sky130_fd_sc_hd__buf_4
Xrepeater689 U$$4244/B2 VGND VGND VPWR VPWR U$$4238/B2 sky130_fd_sc_hd__buf_4
XU$$4371 U$$4508/A1 U$$4381/A2 U$$4510/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4372/A
+ sky130_fd_sc_hd__a22o_1
XU$$4382 U$$4382/A U$$4382/B VGND VGND VPWR VPWR U$$4382/X sky130_fd_sc_hd__xor2_1
XFILLER_65_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4393 U$$4393/A U$$4393/B VGND VGND VPWR VPWR U$$4393/X sky130_fd_sc_hd__xor2_1
XFILLER_77_1137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3670 U$$3805/B1 U$$3566/X U$$3807/B1 U$$3567/X VGND VGND VPWR VPWR U$$3671/A sky130_fd_sc_hd__a22o_1
XU$$3681 U$$3681/A U$$3699/A VGND VGND VPWR VPWR U$$3681/X sky130_fd_sc_hd__xor2_1
XFILLER_77_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3692 U$$4238/B1 U$$3696/A2 U$$4105/A1 U$$3696/B2 VGND VGND VPWR VPWR U$$3693/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_9_0 U$$291/X U$$424/X U$$557/X VGND VGND VPWR VPWR dadda_fa_6_10_0/A dadda_fa_6_9_0/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2980 U$$2980/A U$$3000/B VGND VGND VPWR VPWR U$$2980/X sky130_fd_sc_hd__xor2_1
XU$$2991 U$$2991/A1 U$$2997/A2 U$$2991/B1 U$$2997/B2 VGND VGND VPWR VPWR U$$2992/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_84_2 dadda_fa_4_84_2/A dadda_fa_4_84_2/B dadda_fa_4_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/CIN dadda_fa_5_84_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_77_1 dadda_fa_4_77_1/A dadda_fa_4_77_1/B dadda_fa_4_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/B dadda_fa_5_77_1/B sky130_fd_sc_hd__fa_1
XFILLER_134_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_54_0 dadda_fa_7_54_0/A dadda_fa_7_54_0/B dadda_fa_7_54_0/CIN VGND VGND
+ VPWR VPWR _479_/D _350_/D sky130_fd_sc_hd__fa_1
XFILLER_88_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_670_ _674_/CLK _670_/D VGND VGND VPWR VPWR _670_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$803 U$$938/B1 U$$689/X U$$805/A1 U$$690/X VGND VGND VPWR VPWR U$$804/A sky130_fd_sc_hd__a22o_1
XFILLER_112_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$814 U$$814/A U$$821/A VGND VGND VPWR VPWR U$$814/X sky130_fd_sc_hd__xor2_1
XU$$825 _629_/Q U$$825/B VGND VGND VPWR VPWR U$$825/X sky130_fd_sc_hd__and2_1
XU$$4445_1801 VGND VGND VPWR VPWR U$$4445_1801/HI U$$4445/B sky130_fd_sc_hd__conb_1
XU$$836 U$$973/A1 U$$860/A2 U$$838/A1 U$$860/B2 VGND VGND VPWR VPWR U$$837/A sky130_fd_sc_hd__a22o_1
XFILLER_43_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$847 U$$847/A U$$879/B VGND VGND VPWR VPWR U$$847/X sky130_fd_sc_hd__xor2_1
XFILLER_17_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$858 U$$36/A1 U$$860/A2 U$$38/A1 U$$860/B2 VGND VGND VPWR VPWR U$$859/A sky130_fd_sc_hd__a22o_1
XU$$1008 U$$1008/A U$$980/B VGND VGND VPWR VPWR U$$1008/X sky130_fd_sc_hd__xor2_1
XU$$869 U$$869/A U$$879/B VGND VGND VPWR VPWR U$$869/X sky130_fd_sc_hd__xor2_1
XFILLER_189_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1019 U$$60/A1 U$$1065/A2 U$$62/A1 U$$1065/B2 VGND VGND VPWR VPWR U$$1020/A sky130_fd_sc_hd__a22o_1
XFILLER_32_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_614 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1703 U$$2611/A1 VGND VGND VPWR VPWR U$$8/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_100_clk _634_/CLK VGND VGND VPWR VPWR _495_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_180_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_72_0 dadda_fa_3_72_0/A dadda_fa_3_72_0/B dadda_fa_3_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_0/B dadda_fa_4_72_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_315 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1028 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2210 U$$2895/A1 U$$2248/A2 U$$2210/B1 U$$2248/B2 VGND VGND VPWR VPWR U$$2211/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_34_5 U$$2336/X U$$2366/B input184/X VGND VGND VPWR VPWR dadda_fa_3_35_2/A
+ dadda_fa_4_34_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_101_0 dadda_fa_4_101_0/A dadda_fa_4_101_0/B dadda_fa_4_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/A dadda_fa_5_101_1/A sky130_fd_sc_hd__fa_1
XU$$2221 U$$2221/A U$$2263/B VGND VGND VPWR VPWR U$$2221/X sky130_fd_sc_hd__xor2_1
XU$$2232 U$$449/B1 U$$2248/A2 U$$316/A1 U$$2248/B2 VGND VGND VPWR VPWR U$$2233/A sky130_fd_sc_hd__a22o_1
XU$$2243 U$$2243/A U$$2243/B VGND VGND VPWR VPWR U$$2243/X sky130_fd_sc_hd__xor2_1
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2254 U$$334/B1 U$$2262/A2 U$$201/A1 U$$2262/B2 VGND VGND VPWR VPWR U$$2255/A sky130_fd_sc_hd__a22o_1
XFILLER_90_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2265 U$$2265/A U$$2269/B VGND VGND VPWR VPWR U$$2265/X sky130_fd_sc_hd__xor2_1
XU$$1520 U$$1520/A U$$1558/B VGND VGND VPWR VPWR U$$1520/X sky130_fd_sc_hd__xor2_1
XFILLER_50_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1531 U$$24/A1 U$$1557/A2 U$$985/A1 U$$1557/B2 VGND VGND VPWR VPWR U$$1532/A sky130_fd_sc_hd__a22o_1
XFILLER_90_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2276 U$$3096/B1 U$$2302/A2 U$$3783/B1 U$$2302/B2 VGND VGND VPWR VPWR U$$2277/A
+ sky130_fd_sc_hd__a22o_1
XU$$1542 U$$1542/A U$$1578/B VGND VGND VPWR VPWR U$$1542/X sky130_fd_sc_hd__xor2_1
XU$$2287 U$$2287/A U$$2328/A VGND VGND VPWR VPWR U$$2287/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1553 U$$729/B1 U$$1553/A2 U$$596/A1 U$$1553/B2 VGND VGND VPWR VPWR U$$1554/A sky130_fd_sc_hd__a22o_1
XFILLER_188_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2298 U$$2435/A1 U$$2298/A2 U$$2983/B1 U$$2298/B2 VGND VGND VPWR VPWR U$$2299/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1564 U$$1564/A U$$1588/B VGND VGND VPWR VPWR U$$1564/X sky130_fd_sc_hd__xor2_1
XU$$1575 U$$3354/B1 U$$1577/A2 U$$344/A1 U$$1577/B2 VGND VGND VPWR VPWR U$$1576/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1586 U$$1586/A U$$1588/B VGND VGND VPWR VPWR U$$1586/X sky130_fd_sc_hd__xor2_1
XFILLER_203_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1597 U$$90/A1 U$$1597/A2 U$$92/A1 U$$1597/B2 VGND VGND VPWR VPWR U$$1598/A sky130_fd_sc_hd__a22o_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_94_1 dadda_fa_5_94_1/A dadda_fa_5_94_1/B dadda_fa_5_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_95_0/B dadda_fa_7_94_0/A sky130_fd_sc_hd__fa_1
XFILLER_147_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_87_0 dadda_fa_5_87_0/A dadda_fa_5_87_0/B dadda_fa_5_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_88_0/A dadda_fa_6_87_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_7_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_79_7 U$$3889/X U$$4022/X U$$4155/X VGND VGND VPWR VPWR dadda_fa_2_80_2/CIN
+ dadda_fa_2_79_5/CIN sky130_fd_sc_hd__fa_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$205 final_adder.U$$699/A final_adder.U$$571/B1 final_adder.U$$205/B1
+ VGND VGND VPWR VPWR final_adder.U$$205/X sky130_fd_sc_hd__a21o_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater420 U$$4251/X VGND VGND VPWR VPWR U$$4347/A2 sky130_fd_sc_hd__buf_4
XFILLER_100_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$216 final_adder.U$$711/A final_adder.U$$710/A VGND VGND VPWR VPWR
+ final_adder.U$$300/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$227 final_adder.U$$721/A final_adder.U$$593/B1 final_adder.U$$227/B1
+ VGND VGND VPWR VPWR final_adder.U$$227/X sky130_fd_sc_hd__a21o_1
Xrepeater431 U$$4174/A2 VGND VGND VPWR VPWR U$$4140/A2 sky130_fd_sc_hd__buf_6
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$238 final_adder.U$$733/A final_adder.U$$732/A VGND VGND VPWR VPWR
+ final_adder.U$$310/A sky130_fd_sc_hd__and2_1
XFILLER_211_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater442 U$$98/A2 VGND VGND VPWR VPWR U$$118/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$249 final_adder.U$$743/A final_adder.U$$615/B1 final_adder.U$$249/B1
+ VGND VGND VPWR VPWR final_adder.U$$249/X sky130_fd_sc_hd__a21o_1
Xrepeater453 U$$3977/X VGND VGND VPWR VPWR U$$4107/A2 sky130_fd_sc_hd__buf_4
Xrepeater464 U$$3823/A2 VGND VGND VPWR VPWR U$$3833/A2 sky130_fd_sc_hd__buf_4
Xrepeater475 U$$3664/A2 VGND VGND VPWR VPWR U$$3662/A2 sky130_fd_sc_hd__buf_6
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater486 U$$3418/A2 VGND VGND VPWR VPWR U$$3368/A2 sky130_fd_sc_hd__buf_6
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater497 U$$3283/A2 VGND VGND VPWR VPWR U$$3231/A2 sky130_fd_sc_hd__buf_6
XU$$4190 _588_/Q U$$4196/A2 _589_/Q U$$4196/B2 VGND VGND VPWR VPWR U$$4191/A sky130_fd_sc_hd__a22o_1
XFILLER_129_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4475_1816 VGND VGND VPWR VPWR U$$4475_1816/HI U$$4475/B sky130_fd_sc_hd__conb_1
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_103_2 dadda_fa_3_103_2/A dadda_fa_3_103_2/B dadda_fa_3_103_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_104_1/A dadda_fa_4_103_2/B sky130_fd_sc_hd__fa_1
XFILLER_108_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput201 c[4] VGND VGND VPWR VPWR input201/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_751 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput212 c[5] VGND VGND VPWR VPWR input212/X sky130_fd_sc_hd__clkbuf_4
Xinput223 c[6] VGND VGND VPWR VPWR input223/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput234 c[7] VGND VGND VPWR VPWR input234/X sky130_fd_sc_hd__buf_2
XFILLER_88_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 c[8] VGND VGND VPWR VPWR input245/X sky130_fd_sc_hd__buf_2
XTAP_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput256 c[9] VGND VGND VPWR VPWR input256/X sky130_fd_sc_hd__buf_2
Xdadda_fa_0_67_5 U$$2136/X U$$2269/X U$$2402/X VGND VGND VPWR VPWR dadda_fa_1_68_7/A
+ dadda_fa_2_67_0/A sky130_fd_sc_hd__fa_1
XFILLER_48_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_117_0 dadda_fa_6_117_0/A dadda_fa_6_117_0/B dadda_fa_6_117_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_118_0/B dadda_fa_7_117_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_653_ _662_/CLK _653_/D VGND VGND VPWR VPWR _653_/Q sky130_fd_sc_hd__dfxtp_4
XU$$600 U$$600/A1 U$$600/A2 U$$52/B1 U$$600/B2 VGND VGND VPWR VPWR U$$601/A sky130_fd_sc_hd__a22o_1
XFILLER_91_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$611 U$$611/A U$$613/B VGND VGND VPWR VPWR U$$611/X sky130_fd_sc_hd__xor2_1
XFILLER_112_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_37_3 dadda_fa_3_37_3/A dadda_fa_3_37_3/B dadda_fa_3_37_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_1/B dadda_fa_4_37_2/CIN sky130_fd_sc_hd__fa_1
XU$$622 U$$759/A1 U$$622/A2 U$$624/A1 U$$622/B2 VGND VGND VPWR VPWR U$$623/A sky130_fd_sc_hd__a22o_1
XTAP_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_746 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$633 U$$633/A U$$659/B VGND VGND VPWR VPWR U$$633/X sky130_fd_sc_hd__xor2_1
XU$$644 U$$916/B1 U$$650/A2 U$$781/B1 U$$650/B2 VGND VGND VPWR VPWR U$$645/A sky130_fd_sc_hd__a22o_1
XFILLER_1_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_584_ _588_/CLK _584_/D VGND VGND VPWR VPWR _584_/Q sky130_fd_sc_hd__dfxtp_2
XU$$655 U$$655/A U$$684/A VGND VGND VPWR VPWR U$$655/X sky130_fd_sc_hd__xor2_1
XU$$666 U$$938/B1 U$$668/A2 U$$805/A1 U$$670/B2 VGND VGND VPWR VPWR U$$667/A sky130_fd_sc_hd__a22o_1
XU$$677 U$$677/A U$$685/A VGND VGND VPWR VPWR U$$677/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1015 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$688 U$$810/B U$$688/B VGND VGND VPWR VPWR U$$688/X sky130_fd_sc_hd__and2_1
XFILLER_182_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$699 U$$973/A1 U$$725/A2 U$$838/A1 U$$725/B2 VGND VGND VPWR VPWR U$$700/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_927 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1500 U$$1976/A1 VGND VGND VPWR VPWR U$$880/A1 sky130_fd_sc_hd__buf_6
XFILLER_126_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1511 U$$4027/B1 VGND VGND VPWR VPWR U$$56/A1 sky130_fd_sc_hd__buf_4
Xrepeater1522 U$$4027/A1 VGND VGND VPWR VPWR U$$3342/A1 sky130_fd_sc_hd__buf_4
Xrepeater1533 U$$4160/A1 VGND VGND VPWR VPWR U$$3884/B1 sky130_fd_sc_hd__buf_4
XFILLER_67_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1544 U$$4158/A1 VGND VGND VPWR VPWR U$$2786/B1 sky130_fd_sc_hd__buf_4
Xrepeater1555 _571_/Q VGND VGND VPWR VPWR U$$4154/B1 sky130_fd_sc_hd__buf_6
Xrepeater1566 U$$3876/B1 VGND VGND VPWR VPWR U$$3193/A1 sky130_fd_sc_hd__buf_4
Xrepeater1577 _568_/Q VGND VGND VPWR VPWR U$$4287/A1 sky130_fd_sc_hd__buf_4
Xrepeater1588 U$$856/B1 VGND VGND VPWR VPWR U$$36/A1 sky130_fd_sc_hd__buf_6
XFILLER_125_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1599 U$$3046/B1 VGND VGND VPWR VPWR U$$4007/A1 sky130_fd_sc_hd__buf_6
XFILLER_113_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_32_2 U$$869/X U$$1002/X U$$1135/X VGND VGND VPWR VPWR dadda_fa_3_33_1/A
+ dadda_fa_3_32_3/A sky130_fd_sc_hd__fa_1
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2040 U$$4369/A1 U$$2040/A2 U$$2314/B1 U$$2040/B2 VGND VGND VPWR VPWR U$$2041/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2051 U$$2051/A U$$2054/A VGND VGND VPWR VPWR U$$2051/X sky130_fd_sc_hd__xor2_1
XU$$2062 U$$2062/A U$$2130/B VGND VGND VPWR VPWR U$$2062/X sky130_fd_sc_hd__xor2_1
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2073 U$$2895/A1 U$$2109/A2 U$$2210/B1 U$$2109/B2 VGND VGND VPWR VPWR U$$2074/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2084 U$$2084/A U$$2130/B VGND VGND VPWR VPWR U$$2084/X sky130_fd_sc_hd__xor2_1
XFILLER_210_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1350 U$$1350/A U$$1369/A VGND VGND VPWR VPWR U$$1350/X sky130_fd_sc_hd__xor2_1
XU$$2095 U$$451/A1 U$$2115/A2 U$$999/B1 U$$2115/B2 VGND VGND VPWR VPWR U$$2096/A sky130_fd_sc_hd__a22o_1
XFILLER_211_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1361 U$$948/B1 U$$1367/A2 U$$952/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1362/A sky130_fd_sc_hd__a22o_1
XU$$1372 _637_/Q VGND VGND VPWR VPWR U$$1372/Y sky130_fd_sc_hd__inv_1
XFILLER_22_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1383 U$$1383/A U$$1425/B VGND VGND VPWR VPWR U$$1383/X sky130_fd_sc_hd__xor2_1
XFILLER_188_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1394 U$$435/A1 U$$1424/A2 U$$435/B1 U$$1424/B2 VGND VGND VPWR VPWR U$$1395/A sky130_fd_sc_hd__a22o_1
XFILLER_31_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_692 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_84_5 U$$3367/X U$$3500/X U$$3633/X VGND VGND VPWR VPWR dadda_fa_2_85_3/CIN
+ dadda_fa_2_84_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_77_4 U$$2954/X U$$3087/X U$$3220/X VGND VGND VPWR VPWR dadda_fa_2_78_1/CIN
+ dadda_fa_2_77_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_47_2 dadda_fa_4_47_2/A dadda_fa_4_47_2/B dadda_fa_4_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/CIN dadda_fa_5_47_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_306 _235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_17_0 dadda_fa_7_17_0/A dadda_fa_7_17_0/B dadda_fa_7_17_0/CIN VGND VGND
+ VPWR VPWR _442_/D _313_/D sky130_fd_sc_hd__fa_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_317 _237_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_328 _239_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_339 U$$785/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$90 _514_/Q _386_/Q VGND VGND VPWR VPWR final_adder.U$$585/B1 final_adder.U$$712/A
+ sky130_fd_sc_hd__ha_2
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_832 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_59_3 U$$1322/X U$$1455/X VGND VGND VPWR VPWR dadda_fa_1_60_7/B dadda_fa_2_59_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_122_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1011 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_65_2 U$$935/X U$$1068/X U$$1201/X VGND VGND VPWR VPWR dadda_fa_1_66_6/A
+ dadda_fa_1_65_8/A sky130_fd_sc_hd__fa_1
XFILLER_114_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_42_1 dadda_fa_3_42_1/A dadda_fa_3_42_1/B dadda_fa_3_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_0/CIN dadda_fa_4_42_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_0_58_1 U$$522/X U$$655/X U$$788/X VGND VGND VPWR VPWR dadda_fa_1_59_7/A
+ dadda_fa_1_58_8/B sky130_fd_sc_hd__fa_1
XTAP_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_35_0 dadda_fa_3_35_0/A dadda_fa_3_35_0/B dadda_fa_3_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_0/B dadda_fa_4_35_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$591 final_adder.U$$718/A final_adder.U$$718/B final_adder.U$$591/B1
+ VGND VGND VPWR VPWR final_adder.U$$719/B sky130_fd_sc_hd__a21o_1
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$430 U$$430/A U$$456/B VGND VGND VPWR VPWR U$$430/X sky130_fd_sc_hd__xor2_1
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_636_ _637_/CLK _636_/D VGND VGND VPWR VPWR _636_/Q sky130_fd_sc_hd__dfxtp_1
XU$$441 U$$30/A1 U$$457/A2 U$$32/A1 U$$457/B2 VGND VGND VPWR VPWR U$$442/A sky130_fd_sc_hd__a22o_1
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$452 U$$452/A U$$452/B VGND VGND VPWR VPWR U$$452/X sky130_fd_sc_hd__xor2_1
XFILLER_204_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$463 U$$463/A1 U$$491/A2 U$$463/B1 U$$491/B2 VGND VGND VPWR VPWR U$$464/A sky130_fd_sc_hd__a22o_1
XU$$474 U$$474/A U$$484/B VGND VGND VPWR VPWR U$$474/X sky130_fd_sc_hd__xor2_1
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_567_ _569_/CLK _567_/D VGND VGND VPWR VPWR _567_/Q sky130_fd_sc_hd__dfxtp_2
XU$$485 U$$759/A1 U$$491/A2 U$$624/A1 U$$491/B2 VGND VGND VPWR VPWR U$$486/A sky130_fd_sc_hd__a22o_1
XU$$496 U$$496/A U$$500/B VGND VGND VPWR VPWR U$$496/X sky130_fd_sc_hd__xor2_1
XFILLER_204_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_498_ _500_/CLK _498_/D VGND VGND VPWR VPWR _498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_919 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_94_4 U$$4318/X U$$4451/X input250/X VGND VGND VPWR VPWR dadda_fa_3_95_1/CIN
+ dadda_fa_3_94_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1330 _599_/Q VGND VGND VPWR VPWR U$$4075/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_126_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1341 _597_/Q VGND VGND VPWR VPWR U$$3521/B1 sky130_fd_sc_hd__buf_4
XFILLER_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1352 U$$4480/A1 VGND VGND VPWR VPWR U$$2971/B1 sky130_fd_sc_hd__buf_4
Xrepeater1363 U$$914/A1 VGND VGND VPWR VPWR U$$912/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_87_3 dadda_fa_2_87_3/A dadda_fa_2_87_3/B dadda_fa_2_87_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_1/B dadda_fa_3_87_3/B sky130_fd_sc_hd__fa_1
Xrepeater1374 _593_/Q VGND VGND VPWR VPWR U$$3652/A1 sky130_fd_sc_hd__buf_6
Xrepeater1385 U$$4333/B1 VGND VGND VPWR VPWR U$$4472/A1 sky130_fd_sc_hd__buf_4
Xrepeater1396 U$$3096/B1 VGND VGND VPWR VPWR U$$84/A1 sky130_fd_sc_hd__buf_6
XFILLER_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_57_1 dadda_fa_5_57_1/A dadda_fa_5_57_1/B dadda_fa_5_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_58_0/B dadda_fa_7_57_0/A sky130_fd_sc_hd__fa_2
XFILLER_45_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_103_1 U$$3139/X U$$3272/X U$$3405/X VGND VGND VPWR VPWR dadda_fa_3_104_2/CIN
+ dadda_fa_3_103_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_211_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1180 U$$906/A1 U$$1224/A2 U$$908/A1 U$$1224/B2 VGND VGND VPWR VPWR U$$1181/A sky130_fd_sc_hd__a22o_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1191 U$$1191/A U$$1191/B VGND VGND VPWR VPWR U$$1191/X sky130_fd_sc_hd__xor2_1
XFILLER_52_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_124_0 dadda_fa_5_124_0/A U$$4245/X U$$4378/X VGND VGND VPWR VPWR dadda_fa_6_125_0/B
+ dadda_fa_6_124_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_148_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_982 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_82_2 U$$2033/X U$$2166/X U$$2299/X VGND VGND VPWR VPWR dadda_fa_2_83_2/A
+ dadda_fa_2_82_4/B sky130_fd_sc_hd__fa_1
XFILLER_133_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_75_1 U$$2019/X U$$2152/X U$$2285/X VGND VGND VPWR VPWR dadda_fa_2_76_0/CIN
+ dadda_fa_2_75_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_52_0 dadda_fa_4_52_0/A dadda_fa_4_52_0/B dadda_fa_4_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/A dadda_fa_5_52_1/A sky130_fd_sc_hd__fa_1
XFILLER_58_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_68_0 U$$2537/X U$$2670/X U$$2803/X VGND VGND VPWR VPWR dadda_fa_2_69_0/B
+ dadda_fa_2_68_3/B sky130_fd_sc_hd__fa_1
Xdadda_ha_2_102_3 U$$3802/X U$$3935/X VGND VGND VPWR VPWR dadda_fa_3_103_3/A dadda_fa_4_102_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2809 U$$2809/A U$$2843/B VGND VGND VPWR VPWR U$$2809/X sky130_fd_sc_hd__xor2_1
XANTENNA_103 _287_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_79 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_421_ _627_/CLK _421_/D VGND VGND VPWR VPWR _421_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_136 _290_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _180_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_169 _184_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_clk _628_/CLK VGND VGND VPWR VPWR _648_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _482_/CLK _352_/D VGND VGND VPWR VPWR _352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_283_ _526_/CLK _283_/D VGND VGND VPWR VPWR _283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_97_2 dadda_fa_3_97_2/A dadda_fa_3_97_2/B dadda_fa_3_97_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_1/A dadda_fa_4_97_2/B sky130_fd_sc_hd__fa_1
XFILLER_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_67_0 dadda_fa_6_67_0/A dadda_fa_6_67_0/B dadda_fa_6_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_68_0/B dadda_fa_7_67_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_190_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_70_0 dadda_fa_0_70_0/A U$$546/X U$$679/X VGND VGND VPWR VPWR dadda_fa_1_71_6/B
+ dadda_fa_1_70_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_77_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 a[17] VGND VGND VPWR VPWR _633_/D sky130_fd_sc_hd__clkbuf_2
XTAP_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_119_1 U$$4235/X U$$4368/X U$$4501/X VGND VGND VPWR VPWR dadda_fa_5_120_1/A
+ dadda_fa_5_119_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_5_6_1 U$$418/X U$$452/B VGND VGND VPWR VPWR dadda_fa_6_7_0/B dadda_fa_7_6_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$260 U$$260/A U$$264/B VGND VGND VPWR VPWR U$$260/X sky130_fd_sc_hd__xor2_1
XU$$271 U$$406/B1 U$$141/X U$$271/B1 U$$142/X VGND VGND VPWR VPWR U$$272/A sky130_fd_sc_hd__a22o_1
X_619_ _623_/CLK _619_/D VGND VGND VPWR VPWR _619_/Q sky130_fd_sc_hd__dfxtp_1
XU$$282 U$$8/A1 U$$318/A2 U$$8/B1 U$$318/B2 VGND VGND VPWR VPWR U$$283/A sky130_fd_sc_hd__a22o_1
XFILLER_162_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$293 U$$293/A U$$309/B VGND VGND VPWR VPWR U$$293/X sky130_fd_sc_hd__xor2_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$7 _431_/Q _303_/Q VGND VGND VPWR VPWR final_adder.U$$7/COUT final_adder.U$$7/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_146_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput302 _193_/Q VGND VGND VPWR VPWR o[25] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_1 U$$3383/X U$$3516/X U$$3649/X VGND VGND VPWR VPWR dadda_fa_3_93_0/CIN
+ dadda_fa_3_92_2/CIN sky130_fd_sc_hd__fa_1
Xoutput313 _203_/Q VGND VGND VPWR VPWR o[35] sky130_fd_sc_hd__buf_2
XFILLER_133_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput324 _213_/Q VGND VGND VPWR VPWR o[45] sky130_fd_sc_hd__buf_2
Xoutput335 _223_/Q VGND VGND VPWR VPWR o[55] sky130_fd_sc_hd__buf_2
XFILLER_126_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput346 _233_/Q VGND VGND VPWR VPWR o[65] sky130_fd_sc_hd__buf_2
Xrepeater1160 U$$536/B VGND VGND VPWR VPWR U$$532/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_85_0 U$$3901/X U$$4034/X U$$4167/X VGND VGND VPWR VPWR dadda_fa_3_86_0/B
+ dadda_fa_3_85_2/B sky130_fd_sc_hd__fa_1
XFILLER_114_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1171 U$$411/A VGND VGND VPWR VPWR U$$410/A sky130_fd_sc_hd__buf_6
Xoutput357 _243_/Q VGND VGND VPWR VPWR o[75] sky130_fd_sc_hd__buf_2
Xoutput368 _253_/Q VGND VGND VPWR VPWR o[85] sky130_fd_sc_hd__buf_2
Xrepeater1182 U$$93/B VGND VGND VPWR VPWR U$$57/B sky130_fd_sc_hd__buf_6
Xoutput379 _263_/Q VGND VGND VPWR VPWR o[95] sky130_fd_sc_hd__buf_2
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1193 U$$545/A1 VGND VGND VPWR VPWR U$$4105/B1 sky130_fd_sc_hd__buf_6
XFILLER_141_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_48_7 U$$2896/X U$$3029/X VGND VGND VPWR VPWR dadda_fa_2_49_3/B dadda_fa_3_48_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_7 dadda_fa_1_61_7/A dadda_fa_1_61_7/B dadda_fa_1_61_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_2/CIN dadda_fa_2_61_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_54_6 U$$3174/X U$$3307/X U$$3440/X VGND VGND VPWR VPWR dadda_fa_2_55_2/B
+ dadda_fa_2_54_5/B sky130_fd_sc_hd__fa_1
XFILLER_210_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_47_5 U$$2096/X U$$2229/X U$$2362/X VGND VGND VPWR VPWR dadda_fa_2_48_3/A
+ dadda_fa_2_47_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_167_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_6_0 dadda_fa_7_6_0/A dadda_fa_7_6_0/B dadda_fa_7_6_0/CIN VGND VGND VPWR
+ VPWR _431_/D _302_/D sky130_fd_sc_hd__fa_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_62_clk _535_/CLK VGND VGND VPWR VPWR _582_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_196_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_584 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_84_0 dadda_fa_7_84_0/A dadda_fa_7_84_0/B dadda_fa_7_84_0/CIN VGND VGND
+ VPWR VPWR _509_/D _380_/D sky130_fd_sc_hd__fa_1
XFILLER_13_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4008 U$$4008/A U$$4044/B VGND VGND VPWR VPWR U$$4008/X sky130_fd_sc_hd__xor2_1
XU$$4019 _571_/Q U$$4061/A2 _572_/Q U$$4061/B2 VGND VGND VPWR VPWR U$$4020/A sky130_fd_sc_hd__a22o_1
XFILLER_98_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3307 U$$3307/A U$$3357/B VGND VGND VPWR VPWR U$$3307/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3318 U$$3453/B1 U$$3320/A2 U$$3320/A1 U$$3320/B2 VGND VGND VPWR VPWR U$$3319/A
+ sky130_fd_sc_hd__a22o_1
XU$$3329 U$$3329/A U$$3369/B VGND VGND VPWR VPWR U$$3329/X sky130_fd_sc_hd__xor2_1
XFILLER_24_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2606 U$$2739/A U$$2606/B VGND VGND VPWR VPWR U$$2606/X sky130_fd_sc_hd__and2_1
XFILLER_34_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2617 U$$2754/A1 U$$2663/A2 U$$2756/A1 U$$2663/B2 VGND VGND VPWR VPWR U$$2618/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2628 U$$2628/A U$$2654/B VGND VGND VPWR VPWR U$$2628/X sky130_fd_sc_hd__xor2_1
XU$$2639 U$$2774/B1 U$$2687/A2 U$$2641/A1 U$$2687/B2 VGND VGND VPWR VPWR U$$2640/A
+ sky130_fd_sc_hd__a22o_1
XU$$1905 U$$2314/B1 U$$1909/A2 U$$811/A1 U$$1909/B2 VGND VGND VPWR VPWR U$$1906/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1916 U$$1916/A U$$1916/B VGND VGND VPWR VPWR U$$1916/X sky130_fd_sc_hd__xor2_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1927 U$$1927/A U$$2003/B VGND VGND VPWR VPWR U$$1927/X sky130_fd_sc_hd__xor2_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_53_clk _535_/CLK VGND VGND VPWR VPWR _523_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1938 U$$2210/B1 U$$1976/A2 U$$20/B1 U$$1976/B2 VGND VGND VPWR VPWR U$$1939/A sky130_fd_sc_hd__a22o_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1949 U$$1949/A U$$1957/B VGND VGND VPWR VPWR U$$1949/X sky130_fd_sc_hd__xor2_1
X_404_ _534_/CLK _404_/D VGND VGND VPWR VPWR _404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_335_ _463_/CLK _335_/D VGND VGND VPWR VPWR _335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_266_ _520_/CLK _266_/D VGND VGND VPWR VPWR _266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_197_ _213_/CLK _197_/D VGND VGND VPWR VPWR _197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_64_5 dadda_fa_2_64_5/A dadda_fa_2_64_5/B dadda_fa_2_64_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_2/A dadda_fa_4_64_0/A sky130_fd_sc_hd__fa_2
Xrepeater805 U$$2451/B2 VGND VGND VPWR VPWR U$$2437/B2 sky130_fd_sc_hd__buf_8
XFILLER_116_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater816 U$$2060/X VGND VGND VPWR VPWR U$$2135/B2 sky130_fd_sc_hd__buf_4
XFILLER_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater827 U$$2038/B2 VGND VGND VPWR VPWR U$$2028/B2 sky130_fd_sc_hd__buf_6
Xrepeater838 U$$1786/X VGND VGND VPWR VPWR U$$1907/B2 sky130_fd_sc_hd__buf_8
Xdadda_fa_2_57_4 dadda_fa_2_57_4/A dadda_fa_2_57_4/B dadda_fa_2_57_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/CIN dadda_fa_3_57_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater849 U$$1607/B2 VGND VGND VPWR VPWR U$$1597/B2 sky130_fd_sc_hd__buf_4
XFILLER_37_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$12 U$$12/A1 U$$8/A2 U$$14/A1 U$$8/B2 VGND VGND VPWR VPWR U$$13/A sky130_fd_sc_hd__a22o_1
XU$$23 U$$23/A U$$57/B VGND VGND VPWR VPWR U$$23/X sky130_fd_sc_hd__xor2_1
XU$$34 U$$34/A1 U$$62/A2 U$$36/A1 U$$62/B2 VGND VGND VPWR VPWR U$$35/A sky130_fd_sc_hd__a22o_1
XU$$3830 U$$3830/A U$$3832/B VGND VGND VPWR VPWR U$$3830/X sky130_fd_sc_hd__xor2_1
XU$$3841 U$$3839/B U$$3836/A _672_/Q U$$3836/Y VGND VGND VPWR VPWR U$$3841/X sky130_fd_sc_hd__a22o_4
XU$$45 U$$45/A U$$85/B VGND VGND VPWR VPWR U$$45/X sky130_fd_sc_hd__xor2_1
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$56 U$$56/A1 U$$68/A2 U$$58/A1 U$$68/B2 VGND VGND VPWR VPWR U$$57/A sky130_fd_sc_hd__a22o_1
XU$$67 U$$67/A U$$93/B VGND VGND VPWR VPWR U$$67/X sky130_fd_sc_hd__xor2_1
XU$$3852 U$$4400/A1 U$$3874/A2 _557_/Q U$$3874/B2 VGND VGND VPWR VPWR U$$3853/A sky130_fd_sc_hd__a22o_1
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$78 U$$78/A1 U$$84/A2 U$$80/A1 U$$84/B2 VGND VGND VPWR VPWR U$$79/A sky130_fd_sc_hd__a22o_1
XFILLER_24_107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3863 U$$3863/A U$$3965/B VGND VGND VPWR VPWR U$$3863/X sky130_fd_sc_hd__xor2_1
XU$$3874 U$$584/B1 U$$3874/A2 U$$451/A1 U$$3874/B2 VGND VGND VPWR VPWR U$$3875/A sky130_fd_sc_hd__a22o_1
XU$$3885 U$$3885/A U$$3917/B VGND VGND VPWR VPWR U$$3885/X sky130_fd_sc_hd__xor2_1
XU$$89 U$$89/A U$$93/B VGND VGND VPWR VPWR U$$89/X sky130_fd_sc_hd__xor2_1
XFILLER_52_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3896 U$$4444/A1 U$$3910/A2 U$$3896/B1 U$$3910/B2 VGND VGND VPWR VPWR U$$3897/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_clk _369_/CLK VGND VGND VPWR VPWR _372_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1046 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_14 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_25 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 _282_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_47 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 _285_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_52_3 U$$1574/X U$$1707/X U$$1840/X VGND VGND VPWR VPWR dadda_fa_2_53_1/B
+ dadda_fa_2_52_4/B sky130_fd_sc_hd__fa_1
XFILLER_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_45_2 U$$895/X U$$1028/X U$$1161/X VGND VGND VPWR VPWR dadda_fa_2_46_2/CIN
+ dadda_fa_2_45_5/A sky130_fd_sc_hd__fa_1
XFILLER_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_22_1 dadda_fa_4_22_1/A dadda_fa_4_22_1/B dadda_fa_4_22_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/B dadda_fa_5_22_1/B sky130_fd_sc_hd__fa_1
XFILLER_83_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_38_1 U$$482/X U$$615/X U$$748/X VGND VGND VPWR VPWR dadda_fa_2_39_4/CIN
+ dadda_fa_2_38_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_clk _479_/CLK VGND VGND VPWR VPWR _225_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_4_15_0 U$$303/X U$$436/X U$$569/X VGND VGND VPWR VPWR dadda_fa_5_16_0/A
+ dadda_fa_5_15_1/A sky130_fd_sc_hd__fa_1
XFILLER_19_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_502 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_67_3 dadda_fa_3_67_3/A dadda_fa_3_67_3/B dadda_fa_3_67_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_1/B dadda_fa_4_67_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3104 U$$4474/A1 U$$3148/A2 U$$4476/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3105/A
+ sky130_fd_sc_hd__a22o_1
XU$$3115 U$$3115/A U$$3121/B VGND VGND VPWR VPWR U$$3115/X sky130_fd_sc_hd__xor2_1
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3126 _604_/Q U$$3132/A2 _605_/Q U$$3132/B2 VGND VGND VPWR VPWR U$$3127/A sky130_fd_sc_hd__a22o_1
XU$$3137 U$$3137/A U$$3145/B VGND VGND VPWR VPWR U$$3137/X sky130_fd_sc_hd__xor2_1
XU$$2403 U$$3771/B1 U$$2437/A2 U$$3638/A1 U$$2437/B2 VGND VGND VPWR VPWR U$$2404/A
+ sky130_fd_sc_hd__a22o_1
XU$$3148 U$$3285/A1 U$$3148/A2 U$$3148/B1 U$$3148/B2 VGND VGND VPWR VPWR U$$3149/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2414 U$$2414/A U$$2436/B VGND VGND VPWR VPWR U$$2414/X sky130_fd_sc_hd__xor2_1
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3159 _552_/Q U$$3209/A2 _553_/Q U$$3209/B2 VGND VGND VPWR VPWR U$$3160/A sky130_fd_sc_hd__a22o_1
XU$$2425 U$$3519/B1 U$$2451/A2 U$$3521/B1 U$$2451/B2 VGND VGND VPWR VPWR U$$2426/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2436 U$$2436/A U$$2436/B VGND VGND VPWR VPWR U$$2436/X sky130_fd_sc_hd__xor2_1
XU$$1702 U$$1976/A1 U$$1710/A2 U$$745/A1 U$$1710/B2 VGND VGND VPWR VPWR U$$1703/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2447 U$$392/A1 U$$2451/A2 U$$3132/B1 U$$2451/B2 VGND VGND VPWR VPWR U$$2448/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1713 U$$1713/A U$$1763/B VGND VGND VPWR VPWR U$$1713/X sky130_fd_sc_hd__xor2_1
XU$$2458 U$$2458/A U$$2462/B VGND VGND VPWR VPWR U$$2458/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_26_clk _432_/CLK VGND VGND VPWR VPWR _458_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1724 U$$491/A1 U$$1736/A2 U$$493/A1 U$$1736/B2 VGND VGND VPWR VPWR U$$1725/A sky130_fd_sc_hd__a22o_1
XFILLER_15_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2469 _653_/Q U$$2469/B VGND VGND VPWR VPWR U$$2469/X sky130_fd_sc_hd__and2_1
XFILLER_62_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1735 U$$1735/A U$$1737/B VGND VGND VPWR VPWR U$$1735/X sky130_fd_sc_hd__xor2_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1746 U$$924/A1 U$$1768/A2 U$$924/B1 U$$1768/B2 VGND VGND VPWR VPWR U$$1747/A sky130_fd_sc_hd__a22o_1
XU$$1757 U$$1757/A U$$1763/B VGND VGND VPWR VPWR U$$1757/X sky130_fd_sc_hd__xor2_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1768 U$$946/A1 U$$1768/A2 U$$946/B1 U$$1768/B2 VGND VGND VPWR VPWR U$$1769/A sky130_fd_sc_hd__a22o_1
XFILLER_199_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1779 U$$1779/A U$$1780/A VGND VGND VPWR VPWR U$$1779/X sky130_fd_sc_hd__xor2_1
XFILLER_148_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_318_ _448_/CLK _318_/D VGND VGND VPWR VPWR _318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 a[1] VGND VGND VPWR VPWR _617_/D sky130_fd_sc_hd__clkbuf_2
Xinput23 a[2] VGND VGND VPWR VPWR _618_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 a[3] VGND VGND VPWR VPWR _619_/D sky130_fd_sc_hd__clkbuf_2
X_249_ _253_/CLK _249_/D VGND VGND VPWR VPWR _249_/Q sky130_fd_sc_hd__dfxtp_1
Xinput45 a[4] VGND VGND VPWR VPWR _620_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput56 a[5] VGND VGND VPWR VPWR _621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput67 b[11] VGND VGND VPWR VPWR _563_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput78 b[21] VGND VGND VPWR VPWR _573_/D sky130_fd_sc_hd__clkbuf_1
Xinput89 b[31] VGND VGND VPWR VPWR _583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_782 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_62_2 dadda_fa_2_62_2/A dadda_fa_2_62_2/B dadda_fa_2_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/A dadda_fa_3_62_3/A sky130_fd_sc_hd__fa_1
Xrepeater602 U$$1587/A2 VGND VGND VPWR VPWR U$$1577/A2 sky130_fd_sc_hd__buf_4
XFILLER_96_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater613 U$$259/A2 VGND VGND VPWR VPWR U$$217/A2 sky130_fd_sc_hd__clkbuf_8
Xfinal_adder.U$$409 final_adder.U$$326/B final_adder.U$$646/B final_adder.U$$269/X
+ VGND VGND VPWR VPWR final_adder.U$$650/B sky130_fd_sc_hd__a21o_2
XFILLER_97_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater624 U$$1295/A2 VGND VGND VPWR VPWR U$$1279/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_55_1 dadda_fa_2_55_1/A dadda_fa_2_55_1/B dadda_fa_2_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_0/CIN dadda_fa_3_55_2/CIN sky130_fd_sc_hd__fa_2
Xrepeater635 U$$1194/A2 VGND VGND VPWR VPWR U$$1190/A2 sky130_fd_sc_hd__buf_4
XFILLER_42_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater646 U$$964/X VGND VGND VPWR VPWR U$$1093/B2 sky130_fd_sc_hd__buf_6
Xrepeater657 U$$809/B2 VGND VGND VPWR VPWR U$$765/B2 sky130_fd_sc_hd__buf_4
XFILLER_168_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater668 U$$670/B2 VGND VGND VPWR VPWR U$$622/B2 sky130_fd_sc_hd__buf_4
XU$$4350 U$$4350/A U$$4350/B VGND VGND VPWR VPWR U$$4350/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_32_0 dadda_fa_5_32_0/A dadda_fa_5_32_0/B dadda_fa_5_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_33_0/A dadda_fa_6_32_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_26_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater679 U$$4252/X VGND VGND VPWR VPWR U$$4333/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_48_0 U$$3162/X U$$3295/X U$$3343/B VGND VGND VPWR VPWR dadda_fa_3_49_0/B
+ dadda_fa_3_48_2/B sky130_fd_sc_hd__fa_1
XU$$4361 U$$936/A1 U$$4369/A2 U$$4361/B1 U$$4369/B2 VGND VGND VPWR VPWR U$$4362/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4372 U$$4372/A U$$4383/A VGND VGND VPWR VPWR U$$4372/X sky130_fd_sc_hd__xor2_1
XFILLER_26_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4383 U$$4383/A VGND VGND VPWR VPWR U$$4383/Y sky130_fd_sc_hd__inv_1
XU$$4394 U$$4394/A1 U$$4388/X U$$4396/A1 U$$4438/B2 VGND VGND VPWR VPWR U$$4395/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3660 _597_/Q U$$3664/A2 _598_/Q U$$3664/B2 VGND VGND VPWR VPWR U$$3661/A sky130_fd_sc_hd__a22o_1
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3671 U$$3671/A U$$3671/B VGND VGND VPWR VPWR U$$3671/X sky130_fd_sc_hd__xor2_1
XFILLER_80_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3682 U$$4228/B1 U$$3696/A2 U$$4369/A1 U$$3696/B2 VGND VGND VPWR VPWR U$$3683/A
+ sky130_fd_sc_hd__a22o_1
XU$$3693 U$$3693/A U$$3698/A VGND VGND VPWR VPWR U$$3693/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_17_clk _442_/CLK VGND VGND VPWR VPWR _448_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$2970 U$$2970/A U$$2972/B VGND VGND VPWR VPWR U$$2970/X sky130_fd_sc_hd__xor2_1
XFILLER_179_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_9_1 input256/X dadda_fa_5_9_1/B dadda_ha_4_9_0/SUM VGND VGND VPWR VPWR
+ dadda_fa_6_10_0/B dadda_fa_7_9_0/A sky130_fd_sc_hd__fa_1
XU$$2981 U$$3529/A1 U$$2981/A2 U$$3942/A1 U$$2981/B2 VGND VGND VPWR VPWR U$$2982/A
+ sky130_fd_sc_hd__a22o_1
XU$$2992 U$$2992/A U$$3000/B VGND VGND VPWR VPWR U$$2992/X sky130_fd_sc_hd__xor2_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_502 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_77_2 dadda_fa_4_77_2/A dadda_fa_4_77_2/B dadda_fa_4_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/CIN dadda_fa_5_77_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_47_0 dadda_fa_7_47_0/A dadda_fa_7_47_0/B dadda_fa_7_47_0/CIN VGND VGND
+ VPWR VPWR _472_/D _343_/D sky130_fd_sc_hd__fa_2
XFILLER_130_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_50_0 U$$107/X U$$240/X U$$373/X VGND VGND VPWR VPWR dadda_fa_2_51_0/B
+ dadda_fa_2_50_3/B sky130_fd_sc_hd__fa_1
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$804 U$$804/A U$$804/B VGND VGND VPWR VPWR U$$804/X sky130_fd_sc_hd__xor2_1
XFILLER_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$815 U$$950/B1 U$$819/A2 U$$817/A1 U$$819/B2 VGND VGND VPWR VPWR U$$816/A sky130_fd_sc_hd__a22o_1
XU$$826 U$$824/Y _628_/Q _627_/Q U$$825/X U$$822/Y VGND VGND VPWR VPWR U$$826/X sky130_fd_sc_hd__a32o_4
XFILLER_113_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$837 U$$837/A U$$859/B VGND VGND VPWR VPWR U$$837/X sky130_fd_sc_hd__xor2_1
XFILLER_28_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$848 U$$848/A1 U$$896/A2 U$$848/B1 U$$896/B2 VGND VGND VPWR VPWR U$$849/A sky130_fd_sc_hd__a22o_1
XU$$859 U$$859/A U$$859/B VGND VGND VPWR VPWR U$$859/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1009 U$$48/B1 U$$979/A2 U$$874/A1 U$$979/B2 VGND VGND VPWR VPWR U$$1010/A sky130_fd_sc_hd__a22o_1
XFILLER_83_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1704 U$$2746/B1 VGND VGND VPWR VPWR U$$828/B1 sky130_fd_sc_hd__buf_6
XFILLER_164_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_72_1 dadda_fa_3_72_1/A dadda_fa_3_72_1/B dadda_fa_3_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_0/CIN dadda_fa_4_72_2/A sky130_fd_sc_hd__fa_1
XFILLER_106_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1023 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_65_0 dadda_fa_3_65_0/A dadda_fa_3_65_0/B dadda_fa_3_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_0/B dadda_fa_4_65_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2200 U$$2611/A1 U$$2242/A2 U$$2611/B1 U$$2242/B2 VGND VGND VPWR VPWR U$$2201/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2211 U$$2211/A U$$2243/B VGND VGND VPWR VPWR U$$2211/X sky130_fd_sc_hd__xor2_1
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_101_1 dadda_fa_4_101_1/A dadda_fa_4_101_1/B dadda_fa_4_101_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/B dadda_fa_5_101_1/B sky130_fd_sc_hd__fa_1
XU$$2222 U$$2494/B1 U$$2262/A2 U$$3320/A1 U$$2262/B2 VGND VGND VPWR VPWR U$$2223/A
+ sky130_fd_sc_hd__a22o_1
XU$$2233 U$$2233/A U$$2241/B VGND VGND VPWR VPWR U$$2233/X sky130_fd_sc_hd__xor2_1
XU$$2244 U$$3751/A1 U$$2326/A2 U$$3753/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2245/A
+ sky130_fd_sc_hd__a22o_1
XU$$1510 U$$1642/B U$$1510/B VGND VGND VPWR VPWR U$$1510/X sky130_fd_sc_hd__and2_1
XU$$2255 U$$2255/A U$$2269/B VGND VGND VPWR VPWR U$$2255/X sky130_fd_sc_hd__xor2_1
XU$$1521 U$$2754/A1 U$$1553/A2 U$$2756/A1 U$$1553/B2 VGND VGND VPWR VPWR U$$1522/A
+ sky130_fd_sc_hd__a22o_1
XU$$2266 U$$3771/B1 U$$2274/A2 U$$624/A1 U$$2274/B2 VGND VGND VPWR VPWR U$$2267/A
+ sky130_fd_sc_hd__a22o_1
XU$$1532 U$$1532/A U$$1558/B VGND VGND VPWR VPWR U$$1532/X sky130_fd_sc_hd__xor2_1
XU$$2277 U$$2277/A U$$2303/B VGND VGND VPWR VPWR U$$2277/X sky130_fd_sc_hd__xor2_1
XU$$2288 U$$3519/B1 U$$2326/A2 U$$3521/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2289/A
+ sky130_fd_sc_hd__a22o_1
XU$$1543 U$$582/B1 U$$1561/A2 U$$449/A1 U$$1561/B2 VGND VGND VPWR VPWR U$$1544/A sky130_fd_sc_hd__a22o_1
XFILLER_34_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1554 U$$1554/A U$$1554/B VGND VGND VPWR VPWR U$$1554/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2299 U$$2299/A U$$2299/B VGND VGND VPWR VPWR U$$2299/X sky130_fd_sc_hd__xor2_1
XU$$1565 U$$3346/A1 U$$1587/A2 U$$882/A1 U$$1587/B2 VGND VGND VPWR VPWR U$$1566/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1576 U$$1576/A U$$1578/B VGND VGND VPWR VPWR U$$1576/X sky130_fd_sc_hd__xor2_1
XFILLER_188_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_122_0 dadda_fa_7_122_0/A dadda_fa_7_122_0/B dadda_fa_7_122_0/CIN VGND
+ VGND VPWR VPWR _547_/D _418_/D sky130_fd_sc_hd__fa_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1587 U$$900/B1 U$$1587/A2 U$$82/A1 U$$1587/B2 VGND VGND VPWR VPWR U$$1588/A sky130_fd_sc_hd__a22o_1
XFILLER_176_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1598 U$$1598/A U$$1598/B VGND VGND VPWR VPWR U$$1598/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_87_1 dadda_fa_5_87_1/A dadda_fa_5_87_1/B dadda_fa_5_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_88_0/B dadda_fa_7_87_0/A sky130_fd_sc_hd__fa_2
XFILLER_200_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_6_clk _442_/CLK VGND VGND VPWR VPWR _444_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_171_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_79_8 U$$4288/X U$$4421/X input233/X VGND VGND VPWR VPWR dadda_fa_2_80_3/A
+ dadda_fa_3_79_0/A sky130_fd_sc_hd__fa_2
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$206 final_adder.U$$701/A final_adder.U$$700/A VGND VGND VPWR VPWR
+ final_adder.U$$294/A sky130_fd_sc_hd__and2_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater410 U$$632/A2 VGND VGND VPWR VPWR U$$616/A2 sky130_fd_sc_hd__buf_4
XFILLER_170_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater421 U$$4335/A2 VGND VGND VPWR VPWR U$$4311/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$217 final_adder.U$$711/A final_adder.U$$583/B1 final_adder.U$$217/B1
+ VGND VGND VPWR VPWR final_adder.U$$217/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$228 final_adder.U$$723/A final_adder.U$$722/A VGND VGND VPWR VPWR
+ final_adder.U$$306/B sky130_fd_sc_hd__and2_1
Xrepeater432 U$$4114/X VGND VGND VPWR VPWR U$$4226/A2 sky130_fd_sc_hd__buf_4
Xrepeater443 U$$98/A2 VGND VGND VPWR VPWR U$$84/A2 sky130_fd_sc_hd__buf_4
XFILLER_100_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$239 final_adder.U$$733/A final_adder.U$$605/B1 final_adder.U$$239/B1
+ VGND VGND VPWR VPWR final_adder.U$$239/X sky130_fd_sc_hd__a21o_1
Xrepeater454 U$$3977/X VGND VGND VPWR VPWR U$$4071/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater465 U$$3795/A2 VGND VGND VPWR VPWR U$$3785/A2 sky130_fd_sc_hd__buf_4
XFILLER_84_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater476 U$$3566/X VGND VGND VPWR VPWR U$$3664/A2 sky130_fd_sc_hd__buf_4
XFILLER_211_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater487 U$$3292/X VGND VGND VPWR VPWR U$$3418/A2 sky130_fd_sc_hd__buf_6
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater498 U$$3283/A2 VGND VGND VPWR VPWR U$$3285/A2 sky130_fd_sc_hd__buf_6
XU$$4180 U$$4180/A1 U$$4196/A2 _584_/Q U$$4196/B2 VGND VGND VPWR VPWR U$$4181/A sky130_fd_sc_hd__a22o_1
XFILLER_65_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4191 U$$4191/A U$$4197/B VGND VGND VPWR VPWR U$$4191/X sky130_fd_sc_hd__xor2_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3490 U$$3490/A U$$3490/B VGND VGND VPWR VPWR U$$3490/X sky130_fd_sc_hd__xor2_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_82_0 dadda_fa_4_82_0/A dadda_fa_4_82_0/B dadda_fa_4_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/A dadda_fa_5_82_1/A sky130_fd_sc_hd__fa_1
XFILLER_162_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_103_3 dadda_fa_3_103_3/A dadda_fa_3_103_3/B dadda_fa_3_103_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_104_1/B dadda_fa_4_103_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput202 c[50] VGND VGND VPWR VPWR input202/X sky130_fd_sc_hd__clkbuf_4
Xinput213 c[60] VGND VGND VPWR VPWR input213/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput224 c[70] VGND VGND VPWR VPWR input224/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput235 c[80] VGND VGND VPWR VPWR input235/X sky130_fd_sc_hd__clkbuf_4
XTAP_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput246 c[90] VGND VGND VPWR VPWR input246/X sky130_fd_sc_hd__buf_2
XFILLER_75_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$740 final_adder.U$$740/A final_adder.U$$740/B VGND VGND VPWR VPWR
+ _286_/D sky130_fd_sc_hd__xor2_4
XFILLER_91_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_652_ _662_/CLK _652_/D VGND VGND VPWR VPWR _652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$601 U$$601/A U$$627/B VGND VGND VPWR VPWR U$$601/X sky130_fd_sc_hd__xor2_1
XTAP_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$612 U$$747/B1 U$$616/A2 U$$614/A1 U$$616/B2 VGND VGND VPWR VPWR U$$613/A sky130_fd_sc_hd__a22o_1
XFILLER_1_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$623 U$$623/A U$$665/B VGND VGND VPWR VPWR U$$623/X sky130_fd_sc_hd__xor2_1
XU$$634 U$$84/B1 U$$650/A2 U$$634/B1 U$$650/B2 VGND VGND VPWR VPWR U$$635/A sky130_fd_sc_hd__a22o_1
XU$$645 U$$645/A U$$651/B VGND VGND VPWR VPWR U$$645/X sky130_fd_sc_hd__xor2_1
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_583_ _588_/CLK _583_/D VGND VGND VPWR VPWR _583_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$656 U$$791/B1 U$$682/A2 U$$658/A1 U$$682/B2 VGND VGND VPWR VPWR U$$657/A sky130_fd_sc_hd__a22o_1
XFILLER_204_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$667 U$$667/A U$$669/B VGND VGND VPWR VPWR U$$667/X sky130_fd_sc_hd__xor2_1
XFILLER_17_83 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$678 U$$950/B1 U$$682/A2 U$$678/B1 U$$682/B2 VGND VGND VPWR VPWR U$$679/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$689 U$$687/Y _626_/Q _625_/Q U$$688/X U$$685/Y VGND VGND VPWR VPWR U$$689/X sky130_fd_sc_hd__a32o_4
XFILLER_32_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2189_1730 VGND VGND VPWR VPWR U$$2189_1730/HI U$$2189/B1 sky130_fd_sc_hd__conb_1
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_97_0 dadda_fa_6_97_0/A dadda_fa_6_97_0/B dadda_fa_6_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_98_0/B dadda_fa_7_97_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_200_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1501 U$$3346/A1 VGND VGND VPWR VPWR U$$1976/A1 sky130_fd_sc_hd__buf_4
XFILLER_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1512 U$$4027/B1 VGND VGND VPWR VPWR U$$467/A1 sky130_fd_sc_hd__buf_6
Xrepeater1523 _575_/Q VGND VGND VPWR VPWR U$$4027/A1 sky130_fd_sc_hd__buf_6
Xrepeater1534 U$$50/A1 VGND VGND VPWR VPWR U$$48/B1 sky130_fd_sc_hd__buf_6
XFILLER_4_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1545 U$$4158/A1 VGND VGND VPWR VPWR U$$4432/A1 sky130_fd_sc_hd__buf_8
Xrepeater1556 U$$3741/B1 VGND VGND VPWR VPWR U$$44/A1 sky130_fd_sc_hd__buf_4
XFILLER_4_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1567 U$$3876/B1 VGND VGND VPWR VPWR U$$999/B1 sky130_fd_sc_hd__buf_8
XFILLER_153_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1578 _568_/Q VGND VGND VPWR VPWR U$$3602/A1 sky130_fd_sc_hd__buf_6
Xrepeater1589 U$$719/B1 VGND VGND VPWR VPWR U$$856/B1 sky130_fd_sc_hd__buf_6
XFILLER_154_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_2_33_5 U$$2068/X U$$2201/X VGND VGND VPWR VPWR dadda_fa_3_34_2/A dadda_fa_4_33_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_94_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_32_3 U$$1268/X U$$1401/X U$$1534/X VGND VGND VPWR VPWR dadda_fa_3_33_1/B
+ dadda_fa_3_32_3/B sky130_fd_sc_hd__fa_1
XFILLER_47_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2030 U$$2715/A1 U$$2052/A2 U$$2717/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2031/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2041 U$$2041/A _645_/Q VGND VGND VPWR VPWR U$$2041/X sky130_fd_sc_hd__xor2_1
XU$$2052 U$$2872/B1 U$$2052/A2 U$$2052/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2053/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2063 U$$2746/B1 U$$2129/A2 U$$695/A1 U$$2129/B2 VGND VGND VPWR VPWR U$$2064/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2074 U$$2074/A U$$2108/B VGND VGND VPWR VPWR U$$2074/X sky130_fd_sc_hd__xor2_1
XFILLER_63_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1340 U$$1340/A U$$1369/A VGND VGND VPWR VPWR U$$1340/X sky130_fd_sc_hd__xor2_1
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2085 U$$3453/B1 U$$2129/A2 U$$32/A1 U$$2129/B2 VGND VGND VPWR VPWR U$$2086/A sky130_fd_sc_hd__a22o_1
XU$$1351 U$$253/B1 U$$1367/A2 U$$2721/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1352/A
+ sky130_fd_sc_hd__a22o_1
XU$$2096 U$$2096/A U$$2110/B VGND VGND VPWR VPWR U$$2096/X sky130_fd_sc_hd__xor2_1
XFILLER_210_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1362 U$$1362/A U$$1368/B VGND VGND VPWR VPWR U$$1362/X sky130_fd_sc_hd__xor2_1
XU$$1373 _637_/Q U$$1373/B VGND VGND VPWR VPWR U$$1373/X sky130_fd_sc_hd__and2_1
XFILLER_206_1244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1384 U$$562/A1 U$$1424/A2 U$$973/B1 U$$1424/B2 VGND VGND VPWR VPWR U$$1385/A sky130_fd_sc_hd__a22o_1
XFILLER_200_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1395 U$$1395/A U$$1425/B VGND VGND VPWR VPWR U$$1395/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_77_5 U$$3353/X U$$3486/X U$$3619/X VGND VGND VPWR VPWR dadda_fa_2_78_2/A
+ dadda_fa_2_77_5/A sky130_fd_sc_hd__fa_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_307 _235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_318 _237_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_329 _239_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$80 _504_/Q _376_/Q VGND VGND VPWR VPWR final_adder.U$$575/B1 final_adder.U$$702/A
+ sky130_fd_sc_hd__ha_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$91 _515_/Q _387_/Q VGND VGND VPWR VPWR final_adder.U$$219/B1 final_adder.U$$713/A
+ sky130_fd_sc_hd__ha_2
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1085 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1093_1712 VGND VGND VPWR VPWR U$$1093_1712/HI U$$1093/B1 sky130_fd_sc_hd__conb_1
XFILLER_107_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_101_0 U$$4199/X U$$4332/X U$$4465/X VGND VGND VPWR VPWR dadda_fa_4_102_0/B
+ dadda_fa_4_101_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1023 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_390 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_65_3 U$$1334/X U$$1467/X U$$1600/X VGND VGND VPWR VPWR dadda_fa_1_66_6/B
+ dadda_fa_1_65_8/B sky130_fd_sc_hd__fa_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_42_2 dadda_fa_3_42_2/A dadda_fa_3_42_2/B dadda_fa_3_42_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_1/A dadda_fa_4_42_2/B sky130_fd_sc_hd__fa_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_58_2 U$$921/X U$$1054/X U$$1187/X VGND VGND VPWR VPWR dadda_fa_1_59_7/B
+ dadda_fa_1_58_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_35_1 dadda_fa_3_35_1/A dadda_fa_3_35_1/B dadda_fa_3_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_0/CIN dadda_fa_4_35_2/A sky130_fd_sc_hd__fa_1
XTAP_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$581 final_adder.U$$708/A final_adder.U$$708/B final_adder.U$$581/B1
+ VGND VGND VPWR VPWR final_adder.U$$709/B sky130_fd_sc_hd__a21o_1
XTAP_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_635_ _637_/CLK _635_/D VGND VGND VPWR VPWR _635_/Q sky130_fd_sc_hd__dfxtp_1
XU$$420 U$$420/A U$$452/B VGND VGND VPWR VPWR U$$420/X sky130_fd_sc_hd__xor2_1
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$431 U$$705/A1 U$$457/A2 U$$707/A1 U$$457/B2 VGND VGND VPWR VPWR U$$432/A sky130_fd_sc_hd__a22o_1
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$442 U$$442/A U$$456/B VGND VGND VPWR VPWR U$$442/X sky130_fd_sc_hd__xor2_1
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_12_0 dadda_fa_6_12_0/A dadda_fa_6_12_0/B dadda_fa_6_12_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_13_0/B dadda_fa_7_12_0/CIN sky130_fd_sc_hd__fa_1
XU$$453 U$$999/B1 U$$499/A2 U$$866/A1 U$$499/B2 VGND VGND VPWR VPWR U$$454/A sky130_fd_sc_hd__a22o_1
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_28_0 U$$1526/X U$$1659/X U$$1792/X VGND VGND VPWR VPWR dadda_fa_4_29_0/B
+ dadda_fa_4_28_1/CIN sky130_fd_sc_hd__fa_1
XU$$464 U$$464/A U$$532/B VGND VGND VPWR VPWR U$$464/X sky130_fd_sc_hd__xor2_1
XFILLER_17_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$475 U$$747/B1 U$$483/A2 U$$614/A1 U$$483/B2 VGND VGND VPWR VPWR U$$476/A sky130_fd_sc_hd__a22o_1
X_566_ _566_/CLK _566_/D VGND VGND VPWR VPWR _566_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_588 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$486 U$$486/A U$$536/B VGND VGND VPWR VPWR U$$486/X sky130_fd_sc_hd__xor2_1
XU$$497 U$$84/B1 U$$499/A2 U$$634/B1 U$$499/B2 VGND VGND VPWR VPWR U$$498/A sky130_fd_sc_hd__a22o_1
X_497_ _552_/CLK _497_/D VGND VGND VPWR VPWR _497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1320 U$$3803/A1 VGND VGND VPWR VPWR U$$4214/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_94_5 dadda_fa_2_94_5/A dadda_fa_2_94_5/B dadda_fa_2_94_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_95_2/A dadda_fa_4_94_0/A sky130_fd_sc_hd__fa_1
XFILLER_154_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1331 U$$98/B1 VGND VGND VPWR VPWR U$$648/A1 sky130_fd_sc_hd__buf_4
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1342 U$$918/B1 VGND VGND VPWR VPWR U$$3112/A1 sky130_fd_sc_hd__buf_8
Xrepeater1353 _596_/Q VGND VGND VPWR VPWR U$$4480/A1 sky130_fd_sc_hd__buf_4
Xrepeater1364 U$$3789/B1 VGND VGND VPWR VPWR U$$914/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_87_4 dadda_fa_2_87_4/A dadda_fa_2_87_4/B dadda_fa_2_87_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_1/CIN dadda_fa_3_87_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1375 U$$4474/A1 VGND VGND VPWR VPWR U$$90/A1 sky130_fd_sc_hd__buf_4
XFILLER_141_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1386 _592_/Q VGND VGND VPWR VPWR U$$4333/B1 sky130_fd_sc_hd__buf_6
Xrepeater1397 U$$3783/A1 VGND VGND VPWR VPWR U$$3096/B1 sky130_fd_sc_hd__buf_4
XFILLER_99_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_2_24_1 U$$454/X U$$587/X VGND VGND VPWR VPWR dadda_fa_3_25_3/B dadda_fa_4_24_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_67_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_30_0 U$$67/X U$$200/X U$$333/X VGND VGND VPWR VPWR dadda_fa_3_31_1/A dadda_fa_3_30_2/CIN
+ sky130_fd_sc_hd__fa_2
XFILLER_36_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_103_2 U$$3538/X U$$3671/X U$$3804/X VGND VGND VPWR VPWR dadda_fa_3_104_3/A
+ dadda_fa_4_103_0/A sky130_fd_sc_hd__fa_1
XFILLER_23_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1170 U$$3088/A1 U$$1176/A2 U$$898/A1 U$$1176/B2 VGND VGND VPWR VPWR U$$1171/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1181 U$$1181/A U$$1225/B VGND VGND VPWR VPWR U$$1181/X sky130_fd_sc_hd__xor2_1
XU$$1192 U$$2971/B1 U$$1194/A2 U$$2838/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1193/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_117_0 dadda_fa_5_117_0/A dadda_fa_5_117_0/B dadda_fa_5_117_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_118_0/A dadda_fa_6_117_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_176_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_82_3 U$$2432/X U$$2565/X U$$2698/X VGND VGND VPWR VPWR dadda_fa_2_83_2/B
+ dadda_fa_2_82_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_137_1146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_75_2 U$$2418/X U$$2551/X U$$2684/X VGND VGND VPWR VPWR dadda_fa_2_76_1/A
+ dadda_fa_2_75_4/A sky130_fd_sc_hd__fa_1
XFILLER_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_52_1 dadda_fa_4_52_1/A dadda_fa_4_52_1/B dadda_fa_4_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/B dadda_fa_5_52_1/B sky130_fd_sc_hd__fa_1
XFILLER_59_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_68_1 U$$2936/X U$$3069/X U$$3202/X VGND VGND VPWR VPWR dadda_fa_2_69_0/CIN
+ dadda_fa_2_68_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_45_0 dadda_fa_4_45_0/A dadda_fa_4_45_0/B dadda_fa_4_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/A dadda_fa_5_45_1/A sky130_fd_sc_hd__fa_1
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _287_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_137 _290_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_420_ _626_/CLK _420_/D VGND VGND VPWR VPWR _420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_148 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _180_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_351_ _351_/CLK _351_/D VGND VGND VPWR VPWR _351_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_282_ _526_/CLK _282_/D VGND VGND VPWR VPWR _282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_97_3 dadda_fa_3_97_3/A dadda_fa_3_97_3/B dadda_fa_3_97_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_1/B dadda_fa_4_97_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_496 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_70_1 U$$812/X U$$945/X U$$1078/X VGND VGND VPWR VPWR dadda_fa_1_71_6/CIN
+ dadda_fa_1_70_8/A sky130_fd_sc_hd__fa_1
XTAP_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_0 U$$133/X U$$266/X U$$399/X VGND VGND VPWR VPWR dadda_fa_1_64_5/B
+ dadda_fa_1_63_7/B sky130_fd_sc_hd__fa_1
XTAP_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1066 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$250 U$$250/A U$$250/B VGND VGND VPWR VPWR U$$250/X sky130_fd_sc_hd__xor2_1
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_618_ _633_/CLK _618_/D VGND VGND VPWR VPWR _618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$261 U$$946/A1 U$$263/A2 U$$811/A1 U$$263/B2 VGND VGND VPWR VPWR U$$262/A sky130_fd_sc_hd__a22o_1
XU$$272 U$$272/A U$$272/B VGND VGND VPWR VPWR U$$272/X sky130_fd_sc_hd__xor2_1
XU$$283 U$$283/A U$$319/B VGND VGND VPWR VPWR U$$283/X sky130_fd_sc_hd__xor2_1
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$294 U$$429/B1 U$$308/A2 U$$707/A1 U$$308/B2 VGND VGND VPWR VPWR U$$295/A sky130_fd_sc_hd__a22o_1
XFILLER_162_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_549_ _626_/CLK _549_/D VGND VGND VPWR VPWR _549_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_438 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$0 U$$0/A VGND VGND VPWR VPWR U$$0/Y sky130_fd_sc_hd__inv_1
XFILLER_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$8 _432_/Q _304_/Q VGND VGND VPWR VPWR final_adder.U$$8/COUT final_adder.U$$8/SUM
+ sky130_fd_sc_hd__ha_2
XFILLER_173_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput303 _194_/Q VGND VGND VPWR VPWR o[26] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_2 U$$3782/X U$$3915/X U$$4048/X VGND VGND VPWR VPWR dadda_fa_3_93_1/A
+ dadda_fa_3_92_3/A sky130_fd_sc_hd__fa_1
XFILLER_133_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput314 _204_/Q VGND VGND VPWR VPWR o[36] sky130_fd_sc_hd__buf_2
Xoutput325 _214_/Q VGND VGND VPWR VPWR o[46] sky130_fd_sc_hd__buf_2
Xoutput336 _224_/Q VGND VGND VPWR VPWR o[56] sky130_fd_sc_hd__buf_2
Xrepeater1150 U$$685/A VGND VGND VPWR VPWR U$$684/A sky130_fd_sc_hd__buf_8
Xoutput347 _234_/Q VGND VGND VPWR VPWR o[66] sky130_fd_sc_hd__buf_2
Xrepeater1161 _623_/Q VGND VGND VPWR VPWR U$$536/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_85_1 U$$4300/X U$$4433/X input240/X VGND VGND VPWR VPWR dadda_fa_3_86_0/CIN
+ dadda_fa_3_85_2/CIN sky130_fd_sc_hd__fa_1
Xoutput358 _244_/Q VGND VGND VPWR VPWR o[76] sky130_fd_sc_hd__buf_2
Xrepeater1172 _621_/Q VGND VGND VPWR VPWR U$$411/A sky130_fd_sc_hd__buf_4
Xoutput369 _254_/Q VGND VGND VPWR VPWR o[86] sky130_fd_sc_hd__buf_2
Xrepeater1183 U$$3/A VGND VGND VPWR VPWR U$$93/B sky130_fd_sc_hd__buf_6
Xrepeater1194 U$$817/B1 VGND VGND VPWR VPWR U$$545/A1 sky130_fd_sc_hd__buf_8
XFILLER_82_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_62_0 dadda_fa_5_62_0/A dadda_fa_5_62_0/B dadda_fa_5_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_63_0/A dadda_fa_6_62_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_78_0 dadda_fa_2_78_0/A dadda_fa_2_78_0/B dadda_fa_2_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_0/B dadda_fa_3_78_2/B sky130_fd_sc_hd__fa_1
XFILLER_99_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_8 dadda_fa_1_61_8/A dadda_fa_1_61_8/B dadda_fa_1_61_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_3/A dadda_fa_3_61_0/A sky130_fd_sc_hd__fa_2
XFILLER_45_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_54_7 U$$3573/X U$$3706/X U$$3760/B VGND VGND VPWR VPWR dadda_fa_2_55_2/CIN
+ dadda_fa_2_54_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_894 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_642 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_77_0 dadda_fa_7_77_0/A dadda_fa_7_77_0/B dadda_fa_7_77_0/CIN VGND VGND
+ VPWR VPWR _502_/D _373_/D sky130_fd_sc_hd__fa_1
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_80_0 dadda_fa_1_80_0/A U$$1231/X U$$1364/X VGND VGND VPWR VPWR dadda_fa_2_81_0/CIN
+ dadda_fa_2_80_3/B sky130_fd_sc_hd__fa_1
XFILLER_132_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4009 U$$4418/B1 U$$4065/A2 _567_/Q U$$4065/B2 VGND VGND VPWR VPWR U$$4010/A sky130_fd_sc_hd__a22o_1
XFILLER_59_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3308 U$$3445/A1 U$$3356/A2 U$$3310/A1 U$$3356/B2 VGND VGND VPWR VPWR U$$3309/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3319 U$$3319/A U$$3343/B VGND VGND VPWR VPWR U$$3319/X sky130_fd_sc_hd__xor2_1
XFILLER_207_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_52 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2607 U$$2605/Y _654_/Q U$$2603/A U$$2606/X U$$2603/Y VGND VGND VPWR VPWR U$$2607/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_73_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2618 U$$2618/A U$$2664/B VGND VGND VPWR VPWR U$$2618/X sky130_fd_sc_hd__xor2_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2629 U$$3312/B1 U$$2697/A2 U$$4273/B1 U$$2697/B2 VGND VGND VPWR VPWR U$$2630/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1906 U$$1906/A U$$1916/B VGND VGND VPWR VPWR U$$1906/X sky130_fd_sc_hd__xor2_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1917 U$$1917/A VGND VGND VPWR VPWR U$$1917/Y sky130_fd_sc_hd__inv_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1928 U$$695/A1 U$$1956/A2 U$$2613/B1 U$$1956/B2 VGND VGND VPWR VPWR U$$1929/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1939 U$$1939/A U$$1977/B VGND VGND VPWR VPWR U$$1939/X sky130_fd_sc_hd__xor2_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _559_/CLK _403_/D VGND VGND VPWR VPWR _403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ _463_/CLK _334_/D VGND VGND VPWR VPWR _334_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_265_ _520_/CLK _265_/D VGND VGND VPWR VPWR _265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_196_ _207_/CLK _196_/D VGND VGND VPWR VPWR _196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_95_0 dadda_fa_3_95_0/A dadda_fa_3_95_0/B dadda_fa_3_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_0/B dadda_fa_4_95_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_183_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater806 U$$2334/X VGND VGND VPWR VPWR U$$2451/B2 sky130_fd_sc_hd__buf_6
XFILLER_96_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater817 U$$2115/B2 VGND VGND VPWR VPWR U$$2109/B2 sky130_fd_sc_hd__buf_6
XFILLER_42_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater828 U$$2040/B2 VGND VGND VPWR VPWR U$$2038/B2 sky130_fd_sc_hd__buf_6
Xrepeater839 U$$1736/B2 VGND VGND VPWR VPWR U$$1684/B2 sky130_fd_sc_hd__buf_4
XU$$4510 U$$4510/A1 U$$4388/X U$$4512/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4511/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_57_5 dadda_fa_2_57_5/A dadda_fa_2_57_5/B dadda_fa_2_57_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_2/A dadda_fa_4_57_0/A sky130_fd_sc_hd__fa_2
XU$$13 U$$13/A U$$9/B VGND VGND VPWR VPWR U$$13/X sky130_fd_sc_hd__xor2_1
XFILLER_77_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$24 U$$24/A1 U$$52/A2 U$$26/A1 U$$52/B2 VGND VGND VPWR VPWR U$$25/A sky130_fd_sc_hd__a22o_1
XU$$35 U$$35/A U$$3/A VGND VGND VPWR VPWR U$$35/X sky130_fd_sc_hd__xor2_1
XU$$3820 U$$3820/A U$$3835/A VGND VGND VPWR VPWR U$$3820/X sky130_fd_sc_hd__xor2_1
XU$$3831 U$$406/A1 U$$3833/A2 U$$406/B1 U$$3833/B2 VGND VGND VPWR VPWR U$$3832/A sky130_fd_sc_hd__a22o_1
XU$$46 U$$46/A1 U$$52/A2 U$$48/A1 U$$52/B2 VGND VGND VPWR VPWR U$$47/A sky130_fd_sc_hd__a22o_1
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3842 U$$3842/A1 U$$3874/A2 U$$3844/A1 U$$3874/B2 VGND VGND VPWR VPWR U$$3843/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$57 U$$57/A U$$57/B VGND VGND VPWR VPWR U$$57/X sky130_fd_sc_hd__xor2_1
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3853 U$$3853/A U$$3873/B VGND VGND VPWR VPWR U$$3853/X sky130_fd_sc_hd__xor2_1
XU$$3864 U$$4136/B1 U$$3958/A2 U$$4003/A1 U$$3958/B2 VGND VGND VPWR VPWR U$$3865/A
+ sky130_fd_sc_hd__a22o_1
XU$$68 U$$68/A1 U$$68/A2 U$$70/A1 U$$68/B2 VGND VGND VPWR VPWR U$$69/A sky130_fd_sc_hd__a22o_1
XU$$79 U$$79/A U$$81/B VGND VGND VPWR VPWR U$$79/X sky130_fd_sc_hd__xor2_1
XFILLER_24_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3875 U$$3875/A U$$3895/B VGND VGND VPWR VPWR U$$3875/X sky130_fd_sc_hd__xor2_1
XU$$3886 _573_/Q U$$3916/A2 _574_/Q U$$3916/B2 VGND VGND VPWR VPWR U$$3887/A sky130_fd_sc_hd__a22o_1
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3897 U$$3897/A U$$3933/B VGND VGND VPWR VPWR U$$3897/X sky130_fd_sc_hd__xor2_1
XFILLER_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_15 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_26 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_59 _284_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_931 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_52_4 U$$1973/X U$$2106/X U$$2239/X VGND VGND VPWR VPWR dadda_fa_2_53_1/CIN
+ dadda_fa_2_52_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_56_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_45_3 U$$1294/X U$$1427/X U$$1560/X VGND VGND VPWR VPWR dadda_fa_2_46_3/A
+ dadda_fa_2_45_5/B sky130_fd_sc_hd__fa_1
XFILLER_56_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_22_2 dadda_fa_4_22_2/A dadda_fa_4_22_2/B dadda_fa_4_22_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/CIN dadda_fa_5_22_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_15_1 U$$702/X U$$835/X U$$968/X VGND VGND VPWR VPWR dadda_fa_5_16_0/B
+ dadda_fa_5_15_1/B sky130_fd_sc_hd__fa_1
XFILLER_184_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1027 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_499 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3105 U$$3105/A U$$3107/B VGND VGND VPWR VPWR U$$3105/X sky130_fd_sc_hd__xor2_1
XU$$3116 U$$3799/B1 U$$3120/A2 U$$3529/A1 U$$3120/B2 VGND VGND VPWR VPWR U$$3117/A
+ sky130_fd_sc_hd__a22o_1
XU$$3127 U$$3127/A U$$3133/B VGND VGND VPWR VPWR U$$3127/X sky130_fd_sc_hd__xor2_1
XU$$3138 U$$3412/A1 U$$3144/A2 U$$3412/B1 U$$3144/B2 VGND VGND VPWR VPWR U$$3139/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2404 U$$2404/A U$$2442/B VGND VGND VPWR VPWR U$$2404/X sky130_fd_sc_hd__xor2_1
XU$$3149 U$$3149/A _661_/Q VGND VGND VPWR VPWR U$$3149/X sky130_fd_sc_hd__xor2_1
XU$$2415 U$$2415/A1 U$$2435/A2 U$$3650/A1 U$$2435/B2 VGND VGND VPWR VPWR U$$2416/A
+ sky130_fd_sc_hd__a22o_1
XU$$2426 U$$2426/A U$$2465/A VGND VGND VPWR VPWR U$$2426/X sky130_fd_sc_hd__xor2_1
XFILLER_34_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2437 U$$4490/B1 U$$2437/A2 U$$4357/A1 U$$2437/B2 VGND VGND VPWR VPWR U$$2438/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1703 U$$1703/A U$$1711/B VGND VGND VPWR VPWR U$$1703/X sky130_fd_sc_hd__xor2_1
XU$$2448 U$$2448/A U$$2465/A VGND VGND VPWR VPWR U$$2448/X sky130_fd_sc_hd__xor2_1
XFILLER_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2459 U$$2459/A1 U$$2463/A2 U$$2459/B1 U$$2463/B2 VGND VGND VPWR VPWR U$$2460/A
+ sky130_fd_sc_hd__a22o_1
XU$$1714 U$$3358/A1 U$$1762/A2 U$$2947/B1 U$$1762/B2 VGND VGND VPWR VPWR U$$1715/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1725 U$$1725/A U$$1737/B VGND VGND VPWR VPWR U$$1725/X sky130_fd_sc_hd__xor2_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1736 U$$92/A1 U$$1736/A2 U$$2832/B1 U$$1736/B2 VGND VGND VPWR VPWR U$$1737/A sky130_fd_sc_hd__a22o_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_934 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1747 U$$1747/A U$$1747/B VGND VGND VPWR VPWR U$$1747/X sky130_fd_sc_hd__xor2_1
XU$$1758 U$$2991/A1 U$$1762/A2 U$$2991/B1 U$$1762/B2 VGND VGND VPWR VPWR U$$1759/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1769 U$$1769/A U$$1773/B VGND VGND VPWR VPWR U$$1769/X sky130_fd_sc_hd__xor2_1
XFILLER_202_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_317_ _445_/CLK _317_/D VGND VGND VPWR VPWR _317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 a[20] VGND VGND VPWR VPWR _636_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_248_ _253_/CLK _248_/D VGND VGND VPWR VPWR _248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput24 a[30] VGND VGND VPWR VPWR _646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput35 a[40] VGND VGND VPWR VPWR _656_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput46 a[50] VGND VGND VPWR VPWR _666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput57 a[60] VGND VGND VPWR VPWR _676_/D sky130_fd_sc_hd__clkbuf_1
Xinput68 b[12] VGND VGND VPWR VPWR _564_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_179_ _179_/CLK _179_/D VGND VGND VPWR VPWR _179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput79 b[22] VGND VGND VPWR VPWR _574_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_388 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_62_3 dadda_fa_2_62_3/A dadda_fa_2_62_3/B dadda_fa_2_62_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/B dadda_fa_3_62_3/B sky130_fd_sc_hd__fa_1
XFILLER_97_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater603 U$$1587/A2 VGND VGND VPWR VPWR U$$1561/A2 sky130_fd_sc_hd__buf_4
Xrepeater614 U$$263/A2 VGND VGND VPWR VPWR U$$259/A2 sky130_fd_sc_hd__buf_6
XFILLER_96_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater625 U$$1295/A2 VGND VGND VPWR VPWR U$$1309/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_55_2 dadda_fa_2_55_2/A dadda_fa_2_55_2/B dadda_fa_2_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/A dadda_fa_3_55_3/A sky130_fd_sc_hd__fa_1
Xrepeater636 U$$1208/A2 VGND VGND VPWR VPWR U$$1194/A2 sky130_fd_sc_hd__buf_4
Xrepeater647 U$$964/X VGND VGND VPWR VPWR U$$1065/B2 sky130_fd_sc_hd__buf_6
XFILLER_38_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater658 U$$819/B2 VGND VGND VPWR VPWR U$$783/B2 sky130_fd_sc_hd__buf_4
XFILLER_38_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4340 U$$4340/A U$$4350/B VGND VGND VPWR VPWR U$$4340/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_32_1 dadda_fa_5_32_1/A dadda_fa_5_32_1/B dadda_fa_5_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_33_0/B dadda_fa_7_32_0/A sky130_fd_sc_hd__fa_1
XU$$4351 U$$4351/A1 U$$4381/A2 U$$4353/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4352/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater669 U$$682/B2 VGND VGND VPWR VPWR U$$650/B2 sky130_fd_sc_hd__buf_4
XU$$4362 U$$4362/A U$$4384/A VGND VGND VPWR VPWR U$$4362/X sky130_fd_sc_hd__xor2_1
XFILLER_37_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_48_1 input199/X dadda_fa_2_48_1/B dadda_fa_2_48_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_49_0/CIN dadda_fa_3_48_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_26_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4373 U$$4510/A1 U$$4381/A2 U$$4512/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4374/A
+ sky130_fd_sc_hd__a22o_1
XU$$4384 U$$4384/A VGND VGND VPWR VPWR U$$4384/Y sky130_fd_sc_hd__inv_1
XFILLER_37_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_25_0 dadda_fa_5_25_0/A dadda_fa_5_25_0/B dadda_fa_5_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_26_0/A dadda_fa_6_25_0/CIN sky130_fd_sc_hd__fa_1
XU$$3650 U$$3650/A1 U$$3662/A2 U$$3652/A1 U$$3662/B2 VGND VGND VPWR VPWR U$$3651/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4395 U$$4395/A U$$4395/B VGND VGND VPWR VPWR U$$4395/X sky130_fd_sc_hd__xor2_1
XFILLER_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3661 U$$3661/A U$$3671/B VGND VGND VPWR VPWR U$$3661/X sky130_fd_sc_hd__xor2_1
XU$$3672 U$$3807/B1 U$$3674/A2 U$$4222/A1 U$$3674/B2 VGND VGND VPWR VPWR U$$3673/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3683 U$$3683/A U$$3698/A VGND VGND VPWR VPWR U$$3683/X sky130_fd_sc_hd__xor2_1
XFILLER_80_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3694 U$$4105/A1 U$$3696/A2 U$$4105/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3695/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2960 U$$2960/A U$$2982/B VGND VGND VPWR VPWR U$$2960/X sky130_fd_sc_hd__xor2_1
XU$$2971 U$$4478/A1 U$$2973/A2 U$$2971/B1 U$$2973/B2 VGND VGND VPWR VPWR U$$2972/A
+ sky130_fd_sc_hd__a22o_1
XU$$2982 U$$2982/A U$$2982/B VGND VGND VPWR VPWR U$$2982/X sky130_fd_sc_hd__xor2_1
XU$$2993 _606_/Q U$$2997/A2 _607_/Q U$$2997/B2 VGND VGND VPWR VPWR U$$2994/A sky130_fd_sc_hd__a22o_1
XFILLER_179_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4403_1780 VGND VGND VPWR VPWR U$$4403_1780/HI U$$4403/B sky130_fd_sc_hd__conb_1
XFILLER_147_864 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_1_37_1 U$$480/X U$$613/X VGND VGND VPWR VPWR dadda_fa_2_38_5/A dadda_fa_3_37_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_130_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_50_1 U$$506/X U$$639/X U$$772/X VGND VGND VPWR VPWR dadda_fa_2_51_0/CIN
+ dadda_fa_2_50_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$805 U$$805/A1 U$$689/X U$$805/B1 U$$690/X VGND VGND VPWR VPWR U$$806/A sky130_fd_sc_hd__a22o_1
XFILLER_84_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$816 U$$816/A U$$816/B VGND VGND VPWR VPWR U$$816/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_43_0 U$$93/X U$$226/X U$$359/X VGND VGND VPWR VPWR dadda_fa_2_44_2/CIN
+ dadda_fa_2_43_4/CIN sky130_fd_sc_hd__fa_1
XU$$827 U$$825/B _627_/Q _628_/Q U$$822/Y VGND VGND VPWR VPWR U$$827/X sky130_fd_sc_hd__a22o_4
XU$$838 U$$838/A1 U$$860/A2 U$$840/A1 U$$860/B2 VGND VGND VPWR VPWR U$$839/A sky130_fd_sc_hd__a22o_1
XFILLER_95_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$849 U$$849/A U$$897/B VGND VGND VPWR VPWR U$$849/X sky130_fd_sc_hd__xor2_1
XFILLER_113_76 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_25 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1705 U$$3157/B1 VGND VGND VPWR VPWR U$$967/A1 sky130_fd_sc_hd__buf_4
XFILLER_164_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_72_2 dadda_fa_3_72_2/A dadda_fa_3_72_2/B dadda_fa_3_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_1/A dadda_fa_4_72_2/B sky130_fd_sc_hd__fa_1
XFILLER_117_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_65_1 dadda_fa_3_65_1/A dadda_fa_3_65_1/B dadda_fa_3_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_0/CIN dadda_fa_4_65_2/A sky130_fd_sc_hd__fa_1
XFILLER_152_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_42_0 dadda_fa_6_42_0/A dadda_fa_6_42_0/B dadda_fa_6_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_43_0/B dadda_fa_7_42_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_58_0 dadda_fa_3_58_0/A dadda_fa_3_58_0/B dadda_fa_3_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_0/B dadda_fa_4_58_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_93_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2201 U$$2201/A U$$2241/B VGND VGND VPWR VPWR U$$2201/X sky130_fd_sc_hd__xor2_1
XU$$2212 U$$20/A1 U$$2248/A2 U$$22/A1 U$$2248/B2 VGND VGND VPWR VPWR U$$2213/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_101_2 dadda_fa_4_101_2/A dadda_fa_4_101_2/B dadda_fa_4_101_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/CIN dadda_fa_5_101_1/CIN sky130_fd_sc_hd__fa_1
XU$$2223 U$$2223/A U$$2263/B VGND VGND VPWR VPWR U$$2223/X sky130_fd_sc_hd__xor2_1
XFILLER_62_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2234 U$$2508/A1 U$$2248/A2 U$$2508/B1 U$$2248/B2 VGND VGND VPWR VPWR U$$2235/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2245 U$$2245/A U$$2328/A VGND VGND VPWR VPWR U$$2245/X sky130_fd_sc_hd__xor2_1
XU$$1500 U$$950/B1 U$$1500/A2 U$$817/A1 U$$1500/B2 VGND VGND VPWR VPWR U$$1501/A sky130_fd_sc_hd__a22o_1
XU$$1511 U$$1509/Y _638_/Q U$$1507/A U$$1510/X U$$1507/Y VGND VGND VPWR VPWR U$$1511/X
+ sky130_fd_sc_hd__a32o_2
XU$$2256 U$$201/A1 U$$2262/A2 U$$66/A1 U$$2262/B2 VGND VGND VPWR VPWR U$$2257/A sky130_fd_sc_hd__a22o_1
XU$$2267 U$$2267/A U$$2269/B VGND VGND VPWR VPWR U$$2267/X sky130_fd_sc_hd__xor2_1
XU$$1522 U$$1522/A U$$1554/B VGND VGND VPWR VPWR U$$1522/X sky130_fd_sc_hd__xor2_1
XU$$1533 U$$848/A1 U$$1561/A2 U$$848/B1 U$$1561/B2 VGND VGND VPWR VPWR U$$1534/A sky130_fd_sc_hd__a22o_1
XU$$2278 U$$3783/B1 U$$2298/A2 U$$2963/B1 U$$2298/B2 VGND VGND VPWR VPWR U$$2279/A
+ sky130_fd_sc_hd__a22o_1
XU$$1544 U$$1544/A U$$1562/B VGND VGND VPWR VPWR U$$1544/X sky130_fd_sc_hd__xor2_1
XFILLER_62_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2289 U$$2289/A U$$2328/A VGND VGND VPWR VPWR U$$2289/X sky130_fd_sc_hd__xor2_1
XU$$1555 U$$596/A1 U$$1597/A2 U$$596/B1 U$$1597/B2 VGND VGND VPWR VPWR U$$1556/A sky130_fd_sc_hd__a22o_1
XU$$1566 U$$1566/A U$$1588/B VGND VGND VPWR VPWR U$$1566/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_116_0 dadda_ha_3_116_0/A U$$3697/X VGND VGND VPWR VPWR dadda_fa_4_117_2/CIN
+ dadda_ha_3_116_0/SUM sky130_fd_sc_hd__ha_1
XFILLER_37_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1577 U$$3221/A1 U$$1577/A2 U$$3221/B1 U$$1577/B2 VGND VGND VPWR VPWR U$$1578/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1588 U$$1588/A U$$1588/B VGND VGND VPWR VPWR U$$1588/X sky130_fd_sc_hd__xor2_1
XFILLER_163_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1599 U$$92/A1 U$$1607/A2 U$$2832/B1 U$$1607/B2 VGND VGND VPWR VPWR U$$1600/A sky130_fd_sc_hd__a22o_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_976 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_115_0 dadda_fa_7_115_0/A dadda_fa_7_115_0/B dadda_fa_7_115_0/CIN VGND
+ VGND VPWR VPWR _540_/D _411_/D sky130_fd_sc_hd__fa_1
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_60_0 dadda_fa_2_60_0/A dadda_fa_2_60_0/B dadda_fa_2_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_0/B dadda_fa_3_60_2/B sky130_fd_sc_hd__fa_1
XFILLER_112_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater400 U$$826/X VGND VGND VPWR VPWR U$$948/A2 sky130_fd_sc_hd__buf_8
XU$$4433_1795 VGND VGND VPWR VPWR U$$4433_1795/HI U$$4433/B sky130_fd_sc_hd__conb_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$207 final_adder.U$$701/A final_adder.U$$573/B1 final_adder.U$$207/B1
+ VGND VGND VPWR VPWR final_adder.U$$207/X sky130_fd_sc_hd__a21o_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater411 U$$632/A2 VGND VGND VPWR VPWR U$$600/A2 sky130_fd_sc_hd__buf_8
XFILLER_111_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater422 U$$4335/A2 VGND VGND VPWR VPWR U$$4327/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_85_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$218 final_adder.U$$713/A final_adder.U$$712/A VGND VGND VPWR VPWR
+ final_adder.U$$300/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$229 final_adder.U$$723/A final_adder.U$$595/B1 final_adder.U$$229/B1
+ VGND VGND VPWR VPWR final_adder.U$$229/X sky130_fd_sc_hd__a21o_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater433 U$$4244/A2 VGND VGND VPWR VPWR U$$4238/A2 sky130_fd_sc_hd__buf_4
XFILLER_85_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater444 U$$98/A2 VGND VGND VPWR VPWR U$$128/A2 sky130_fd_sc_hd__buf_4
Xrepeater455 U$$3932/A2 VGND VGND VPWR VPWR U$$3916/A2 sky130_fd_sc_hd__buf_4
Xrepeater466 U$$3805/A2 VGND VGND VPWR VPWR U$$3795/A2 sky130_fd_sc_hd__buf_4
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater477 U$$3566/X VGND VGND VPWR VPWR U$$3674/A2 sky130_fd_sc_hd__buf_6
XU$$4170 U$$4444/A1 U$$4226/A2 U$$4444/B1 U$$4226/B2 VGND VGND VPWR VPWR U$$4171/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater488 U$$3378/A2 VGND VGND VPWR VPWR U$$3320/A2 sky130_fd_sc_hd__buf_6
XU$$4181 U$$4181/A U$$4197/B VGND VGND VPWR VPWR U$$4181/X sky130_fd_sc_hd__xor2_1
Xrepeater499 U$$3273/A2 VGND VGND VPWR VPWR U$$3263/A2 sky130_fd_sc_hd__buf_4
XU$$4509_1833 VGND VGND VPWR VPWR U$$4509_1833/HI U$$4509/B sky130_fd_sc_hd__conb_1
XU$$4192 _589_/Q U$$4196/A2 _590_/Q U$$4196/B2 VGND VGND VPWR VPWR U$$4193/A sky130_fd_sc_hd__a22o_1
XFILLER_93_692 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3480 U$$3480/A U$$3490/B VGND VGND VPWR VPWR U$$3480/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3491 U$$3626/B1 U$$3537/A2 U$$4450/B1 U$$3537/B2 VGND VGND VPWR VPWR U$$3492/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2790 U$$596/B1 U$$2798/A2 U$$463/A1 U$$2798/B2 VGND VGND VPWR VPWR U$$2791/A sky130_fd_sc_hd__a22o_1
XFILLER_43_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_82_1 dadda_fa_4_82_1/A dadda_fa_4_82_1/B dadda_fa_4_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/B dadda_fa_5_82_1/B sky130_fd_sc_hd__fa_1
XFILLER_135_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_75_0 dadda_fa_4_75_0/A dadda_fa_4_75_0/B dadda_fa_4_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/A dadda_fa_5_75_1/A sky130_fd_sc_hd__fa_1
XFILLER_134_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput203 c[51] VGND VGND VPWR VPWR input203/X sky130_fd_sc_hd__clkbuf_4
Xinput214 c[61] VGND VGND VPWR VPWR input214/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput225 c[71] VGND VGND VPWR VPWR input225/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput236 c[81] VGND VGND VPWR VPWR input236/X sky130_fd_sc_hd__clkbuf_4
XFILLER_75_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput247 c[91] VGND VGND VPWR VPWR input247/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$730 final_adder.U$$730/A final_adder.U$$730/B VGND VGND VPWR VPWR
+ _276_/D sky130_fd_sc_hd__xor2_4
XTAP_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$741 final_adder.U$$741/A final_adder.U$$741/B VGND VGND VPWR VPWR
+ _287_/D sky130_fd_sc_hd__xor2_4
X_651_ _662_/CLK _651_/D VGND VGND VPWR VPWR _651_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$602 U$$876/A1 U$$616/A2 U$$878/A1 U$$616/B2 VGND VGND VPWR VPWR U$$603/A sky130_fd_sc_hd__a22o_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$613 U$$613/A U$$613/B VGND VGND VPWR VPWR U$$613/X sky130_fd_sc_hd__xor2_1
XFILLER_29_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$624 U$$624/A1 U$$632/A2 U$$624/B1 U$$632/B2 VGND VGND VPWR VPWR U$$625/A sky130_fd_sc_hd__a22o_1
X_582_ _582_/CLK _582_/D VGND VGND VPWR VPWR _582_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$635 U$$635/A U$$651/B VGND VGND VPWR VPWR U$$635/X sky130_fd_sc_hd__xor2_1
XU$$646 U$$781/B1 U$$650/A2 U$$648/A1 U$$650/B2 VGND VGND VPWR VPWR U$$647/A sky130_fd_sc_hd__a22o_1
XFILLER_71_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$657 U$$657/A U$$684/A VGND VGND VPWR VPWR U$$657/X sky130_fd_sc_hd__xor2_1
XFILLER_189_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$668 U$$805/A1 U$$668/A2 U$$805/B1 U$$670/B2 VGND VGND VPWR VPWR U$$669/A sky130_fd_sc_hd__a22o_1
XFILLER_71_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$679 U$$679/A U$$684/A VGND VGND VPWR VPWR U$$679/X sky130_fd_sc_hd__xor2_1
XFILLER_72_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1502 U$$2796/B1 VGND VGND VPWR VPWR U$$58/A1 sky130_fd_sc_hd__buf_4
Xrepeater1513 U$$4440/A1 VGND VGND VPWR VPWR U$$4301/B1 sky130_fd_sc_hd__buf_4
XFILLER_32_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1524 _574_/Q VGND VGND VPWR VPWR U$$4436/A1 sky130_fd_sc_hd__buf_4
XFILLER_181_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1535 U$$733/B1 VGND VGND VPWR VPWR U$$596/B1 sky130_fd_sc_hd__buf_6
Xrepeater1546 _572_/Q VGND VGND VPWR VPWR U$$4158/A1 sky130_fd_sc_hd__buf_6
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1557 U$$3056/B1 VGND VGND VPWR VPWR U$$42/B1 sky130_fd_sc_hd__buf_4
Xrepeater1568 U$$4426/A1 VGND VGND VPWR VPWR U$$3876/B1 sky130_fd_sc_hd__buf_6
XFILLER_4_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1579 U$$584/B1 VGND VGND VPWR VPWR U$$449/A1 sky130_fd_sc_hd__buf_6
XFILLER_154_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2020 U$$3388/B1 U$$2028/A2 U$$3253/B1 U$$2028/B2 VGND VGND VPWR VPWR U$$2021/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_32_4 U$$1667/X U$$1800/X U$$1933/X VGND VGND VPWR VPWR dadda_fa_3_33_1/CIN
+ dadda_fa_3_32_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2031 U$$2031/A U$$2054/A VGND VGND VPWR VPWR U$$2031/X sky130_fd_sc_hd__xor2_1
XFILLER_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2042 U$$2314/B1 U$$2052/A2 U$$946/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2043/A
+ sky130_fd_sc_hd__a22o_1
XU$$2053 U$$2053/A U$$2054/A VGND VGND VPWR VPWR U$$2053/X sky130_fd_sc_hd__xor2_1
XFILLER_50_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2064 U$$2064/A U$$2130/B VGND VGND VPWR VPWR U$$2064/X sky130_fd_sc_hd__xor2_1
XU$$2075 U$$2210/B1 U$$2115/A2 U$$20/B1 U$$2115/B2 VGND VGND VPWR VPWR U$$2076/A sky130_fd_sc_hd__a22o_1
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1330 U$$1330/A U$$1332/B VGND VGND VPWR VPWR U$$1330/X sky130_fd_sc_hd__xor2_1
XU$$2086 U$$2086/A U$$2130/B VGND VGND VPWR VPWR U$$2086/X sky130_fd_sc_hd__xor2_1
XU$$1341 U$$791/B1 U$$1345/A2 U$$4357/A1 U$$1345/B2 VGND VGND VPWR VPWR U$$1342/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1352 U$$1352/A U$$1368/B VGND VGND VPWR VPWR U$$1352/X sky130_fd_sc_hd__xor2_1
XU$$2097 U$$316/A1 U$$2109/A2 U$$3741/B1 U$$2109/B2 VGND VGND VPWR VPWR U$$2098/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1363 U$$950/B1 U$$1367/A2 U$$817/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1364/A sky130_fd_sc_hd__a22o_1
XFILLER_50_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1374 U$$1372/Y _636_/Q U$$1370/A U$$1373/X U$$1370/Y VGND VGND VPWR VPWR U$$1374/X
+ sky130_fd_sc_hd__a32o_4
XU$$1385 U$$1385/A U$$1425/B VGND VGND VPWR VPWR U$$1385/X sky130_fd_sc_hd__xor2_1
XFILLER_206_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1396 U$$435/B1 U$$1424/A2 U$$302/A1 U$$1424/B2 VGND VGND VPWR VPWR U$$1397/A sky130_fd_sc_hd__a22o_1
XFILLER_200_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_106_0_1865 VGND VGND VPWR VPWR dadda_fa_2_106_0/A dadda_fa_2_106_0_1865/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_135_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_92_0 dadda_fa_5_92_0/A dadda_fa_5_92_0/B dadda_fa_5_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_93_0/A dadda_fa_6_92_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_190_214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_77_6 U$$3752/X U$$3885/X U$$4018/X VGND VGND VPWR VPWR dadda_fa_2_78_2/B
+ dadda_fa_2_77_5/B sky130_fd_sc_hd__fa_1
XFILLER_86_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 _235_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_319 _237_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$70 _494_/Q _366_/Q VGND VGND VPWR VPWR final_adder.U$$565/B1 final_adder.U$$692/A
+ sky130_fd_sc_hd__ha_2
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$81 _505_/Q _377_/Q VGND VGND VPWR VPWR final_adder.U$$209/B1 final_adder.U$$703/A
+ sky130_fd_sc_hd__ha_1
XFILLER_110_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$92 _516_/Q _388_/Q VGND VGND VPWR VPWR final_adder.U$$587/B1 final_adder.U$$714/A
+ sky130_fd_sc_hd__ha_1
XFILLER_80_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1097 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_101_1 input131/X dadda_fa_3_101_1/B dadda_fa_3_101_1/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_102_0/CIN dadda_fa_4_101_2/A sky130_fd_sc_hd__fa_1
XFILLER_102_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_122_0 dadda_fa_6_122_0/A dadda_fa_6_122_0/B dadda_fa_6_122_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_123_0/B dadda_fa_7_122_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_65_4 U$$1733/X U$$1866/X U$$1999/X VGND VGND VPWR VPWR dadda_fa_1_66_6/CIN
+ dadda_fa_1_65_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_42_3 dadda_fa_3_42_3/A dadda_fa_3_42_3/B dadda_fa_3_42_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_1/B dadda_fa_4_42_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_36_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$571 final_adder.U$$698/A final_adder.U$$698/B final_adder.U$$571/B1
+ VGND VGND VPWR VPWR final_adder.U$$699/B sky130_fd_sc_hd__a21o_1
XTAP_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_634_ _634_/CLK _634_/D VGND VGND VPWR VPWR _634_/Q sky130_fd_sc_hd__dfxtp_1
XU$$410 U$$410/A VGND VGND VPWR VPWR U$$410/Y sky130_fd_sc_hd__inv_1
XTAP_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_35_2 dadda_fa_3_35_2/A dadda_fa_3_35_2/B dadda_fa_3_35_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_1/A dadda_fa_4_35_2/B sky130_fd_sc_hd__fa_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$421 U$$556/B1 U$$447/A2 U$$695/B1 U$$447/B2 VGND VGND VPWR VPWR U$$422/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$593 final_adder.U$$720/A final_adder.U$$720/B final_adder.U$$593/B1
+ VGND VGND VPWR VPWR final_adder.U$$721/B sky130_fd_sc_hd__a21o_1
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$432 U$$432/A U$$456/B VGND VGND VPWR VPWR U$$432/X sky130_fd_sc_hd__xor2_1
XFILLER_205_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$443 U$$715/B1 U$$447/A2 U$$582/A1 U$$447/B2 VGND VGND VPWR VPWR U$$444/A sky130_fd_sc_hd__a22o_1
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$454 U$$454/A U$$500/B VGND VGND VPWR VPWR U$$454/X sky130_fd_sc_hd__xor2_1
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_565_ _569_/CLK _565_/D VGND VGND VPWR VPWR _565_/Q sky130_fd_sc_hd__dfxtp_4
Xdadda_fa_3_28_1 U$$1925/X U$$2003/B input177/X VGND VGND VPWR VPWR dadda_fa_4_29_0/CIN
+ dadda_fa_4_28_2/A sky130_fd_sc_hd__fa_1
XFILLER_45_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$465 U$$54/A1 U$$499/A2 U$$56/A1 U$$499/B2 VGND VGND VPWR VPWR U$$466/A sky130_fd_sc_hd__a22o_1
XU$$476 U$$476/A U$$484/B VGND VGND VPWR VPWR U$$476/X sky130_fd_sc_hd__xor2_1
XFILLER_45_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$487 U$$624/A1 U$$415/X U$$624/B1 U$$416/X VGND VGND VPWR VPWR U$$488/A sky130_fd_sc_hd__a22o_1
XFILLER_32_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$498 U$$498/A U$$500/B VGND VGND VPWR VPWR U$$498/X sky130_fd_sc_hd__xor2_1
X_496_ _496_/CLK _496_/D VGND VGND VPWR VPWR _496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1310 U$$4353/A1 VGND VGND VPWR VPWR U$$928/A1 sky130_fd_sc_hd__buf_6
Xrepeater1321 U$$3529/A1 VGND VGND VPWR VPWR U$$3803/A1 sky130_fd_sc_hd__buf_4
Xrepeater1332 U$$3386/B1 VGND VGND VPWR VPWR U$$98/B1 sky130_fd_sc_hd__buf_6
Xrepeater1343 U$$4482/A1 VGND VGND VPWR VPWR U$$2838/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1354 _596_/Q VGND VGND VPWR VPWR U$$3658/A1 sky130_fd_sc_hd__buf_6
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_526 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_87_5 dadda_fa_2_87_5/A dadda_fa_2_87_5/B dadda_fa_2_87_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_2/A dadda_fa_4_87_0/A sky130_fd_sc_hd__fa_1
Xrepeater1365 U$$3380/A1 VGND VGND VPWR VPWR U$$229/A1 sky130_fd_sc_hd__buf_8
XFILLER_158_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1376 U$$4472/B1 VGND VGND VPWR VPWR U$$4474/A1 sky130_fd_sc_hd__clkbuf_8
Xrepeater1387 U$$4194/B1 VGND VGND VPWR VPWR U$$908/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_125_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1398 U$$4468/A1 VGND VGND VPWR VPWR U$$3783/A1 sky130_fd_sc_hd__buf_4
XFILLER_141_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_30_1 U$$466/X U$$599/X U$$732/X VGND VGND VPWR VPWR dadda_fa_3_31_1/B
+ dadda_fa_3_30_3/A sky130_fd_sc_hd__fa_1
XFILLER_169_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1018 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1160 U$$201/A1 U$$1190/A2 U$$749/B1 U$$1190/B2 VGND VGND VPWR VPWR U$$1161/A sky130_fd_sc_hd__a22o_1
XFILLER_195_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1171 U$$1171/A U$$1177/B VGND VGND VPWR VPWR U$$1171/X sky130_fd_sc_hd__xor2_1
XU$$1182 U$$2415/A1 U$$1224/A2 U$$3650/A1 U$$1224/B2 VGND VGND VPWR VPWR U$$1183/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1193 U$$1193/A U$$1203/B VGND VGND VPWR VPWR U$$1193/X sky130_fd_sc_hd__xor2_1
XFILLER_148_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_117_1 dadda_fa_5_117_1/A dadda_fa_5_117_1/B dadda_fa_5_117_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_118_0/B dadda_fa_7_117_0/A sky130_fd_sc_hd__fa_1
XFILLER_40_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_439 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_578 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_494 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_82_4 U$$2831/X U$$2964/X U$$3097/X VGND VGND VPWR VPWR dadda_fa_2_83_2/CIN
+ dadda_fa_2_82_5/A sky130_fd_sc_hd__fa_1
XFILLER_172_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_75_3 U$$2817/X U$$2950/X U$$3083/X VGND VGND VPWR VPWR dadda_fa_2_76_1/B
+ dadda_fa_2_75_4/B sky130_fd_sc_hd__fa_1
XFILLER_160_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_52_2 dadda_fa_4_52_2/A dadda_fa_4_52_2/B dadda_fa_4_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/CIN dadda_fa_5_52_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_131_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_2 U$$3335/X U$$3468/X U$$3601/X VGND VGND VPWR VPWR dadda_fa_2_69_1/A
+ dadda_fa_2_68_4/A sky130_fd_sc_hd__fa_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_45_1 dadda_fa_4_45_1/A dadda_fa_4_45_1/B dadda_fa_4_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/B dadda_fa_5_45_1/B sky130_fd_sc_hd__fa_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_22_0 dadda_fa_7_22_0/A dadda_fa_7_22_0/B dadda_fa_7_22_0/CIN VGND VGND
+ VPWR VPWR _447_/D _318_/D sky130_fd_sc_hd__fa_1
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_0 dadda_fa_4_38_0/A dadda_fa_4_38_0/B dadda_fa_4_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/A dadda_fa_5_38_1/A sky130_fd_sc_hd__fa_1
XFILLER_27_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _287_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_138 _290_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_350_ _351_/CLK _350_/D VGND VGND VPWR VPWR _350_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_281_ _526_/CLK _281_/D VGND VGND VPWR VPWR _281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_807 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_57_2 U$$919/X U$$1052/X VGND VGND VPWR VPWR dadda_fa_1_58_7/CIN dadda_fa_2_57_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_70_2 U$$1211/X U$$1344/X U$$1477/X VGND VGND VPWR VPWR dadda_fa_1_71_7/A
+ dadda_fa_1_70_8/B sky130_fd_sc_hd__fa_1
XFILLER_104_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_1 U$$532/X U$$665/X U$$798/X VGND VGND VPWR VPWR dadda_fa_1_64_5/CIN
+ dadda_fa_1_63_7/CIN sky130_fd_sc_hd__fa_1
XTAP_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_40_0 dadda_fa_3_40_0/A dadda_fa_3_40_0/B dadda_fa_3_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_0/B dadda_fa_4_40_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_56_0 U$$119/X U$$252/X U$$385/X VGND VGND VPWR VPWR dadda_fa_1_57_7/B
+ dadda_fa_1_56_8/B sky130_fd_sc_hd__fa_1
XFILLER_65_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$240 U$$240/A U$$250/B VGND VGND VPWR VPWR U$$240/X sky130_fd_sc_hd__xor2_1
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$251 U$$251/A1 U$$259/A2 U$$251/B1 U$$259/B2 VGND VGND VPWR VPWR U$$252/A sky130_fd_sc_hd__a22o_1
X_617_ _623_/CLK _617_/D VGND VGND VPWR VPWR _617_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$262 U$$262/A U$$264/B VGND VGND VPWR VPWR U$$262/X sky130_fd_sc_hd__xor2_1
XFILLER_91_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$273 _619_/Q VGND VGND VPWR VPWR U$$273/Y sky130_fd_sc_hd__inv_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$284 U$$8/B1 U$$318/A2 U$$12/A1 U$$318/B2 VGND VGND VPWR VPWR U$$285/A sky130_fd_sc_hd__a22o_1
XFILLER_60_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_548_ _626_/CLK _548_/D VGND VGND VPWR VPWR _548_/Q sky130_fd_sc_hd__dfxtp_1
XU$$295 U$$295/A U$$309/B VGND VGND VPWR VPWR U$$295/X sky130_fd_sc_hd__xor2_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_479_ _479_/CLK _479_/D VGND VGND VPWR VPWR _479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1095 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1 U$$1/A VGND VGND VPWR VPWR U$$3/B sky130_fd_sc_hd__inv_1
XFILLER_127_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$9 _433_/Q _305_/Q VGND VGND VPWR VPWR final_adder.U$$9/COUT final_adder.U$$9/SUM
+ sky130_fd_sc_hd__ha_2
XFILLER_145_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput304 _195_/Q VGND VGND VPWR VPWR o[27] sky130_fd_sc_hd__buf_2
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_92_3 U$$4181/X U$$4314/X U$$4447/X VGND VGND VPWR VPWR dadda_fa_3_93_1/B
+ dadda_fa_3_92_3/B sky130_fd_sc_hd__fa_1
Xoutput315 _205_/Q VGND VGND VPWR VPWR o[37] sky130_fd_sc_hd__buf_2
XFILLER_114_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput326 _215_/Q VGND VGND VPWR VPWR o[47] sky130_fd_sc_hd__buf_2
XFILLER_126_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1140 U$$804/B VGND VGND VPWR VPWR U$$796/B sky130_fd_sc_hd__buf_6
Xoutput337 _225_/Q VGND VGND VPWR VPWR o[57] sky130_fd_sc_hd__buf_2
Xrepeater1151 U$$669/B VGND VGND VPWR VPWR U$$589/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_85_2 dadda_fa_2_85_2/A dadda_fa_2_85_2/B dadda_fa_2_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/A dadda_fa_3_85_3/A sky130_fd_sc_hd__fa_1
Xrepeater1162 U$$547/A VGND VGND VPWR VPWR U$$518/B sky130_fd_sc_hd__buf_6
Xoutput348 _235_/Q VGND VGND VPWR VPWR o[67] sky130_fd_sc_hd__buf_2
XFILLER_82_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput359 _245_/Q VGND VGND VPWR VPWR o[77] sky130_fd_sc_hd__buf_2
Xrepeater1173 U$$226/B VGND VGND VPWR VPWR U$$190/B sky130_fd_sc_hd__buf_6
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1184 U$$2/A VGND VGND VPWR VPWR U$$3/A sky130_fd_sc_hd__buf_4
Xrepeater1195 U$$2872/B1 VGND VGND VPWR VPWR U$$817/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_5_62_1 dadda_fa_5_62_1/A dadda_fa_5_62_1/B dadda_fa_5_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_63_0/B dadda_fa_7_62_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_78_1 dadda_fa_2_78_1/A dadda_fa_2_78_1/B dadda_fa_2_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_0/CIN dadda_fa_3_78_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_54 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_55_0 dadda_fa_5_55_0/A dadda_fa_5_55_0/B dadda_fa_5_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_56_0/A dadda_fa_6_55_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_8 input206/X dadda_fa_1_54_8/B dadda_fa_1_54_8/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_55_3/A dadda_fa_3_54_0/A sky130_fd_sc_hd__fa_2
XFILLER_209_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_101_0 U$$2602/Y U$$2736/X U$$2869/X VGND VGND VPWR VPWR dadda_fa_3_102_1/CIN
+ dadda_fa_3_101_3/A sky130_fd_sc_hd__fa_1
XFILLER_36_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_80_1 U$$1497/X U$$1630/X U$$1763/X VGND VGND VPWR VPWR dadda_fa_2_81_1/A
+ dadda_fa_2_80_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_73_0 U$$1882/X U$$2015/X U$$2148/X VGND VGND VPWR VPWR dadda_fa_2_74_0/B
+ dadda_fa_2_73_3/B sky130_fd_sc_hd__fa_1
XFILLER_63_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3309 U$$3309/A U$$3357/B VGND VGND VPWR VPWR U$$3309/X sky130_fd_sc_hd__xor2_1
XFILLER_86_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2608 U$$2606/B U$$2603/A _654_/Q U$$2603/Y VGND VGND VPWR VPWR U$$2608/X sky130_fd_sc_hd__a22o_4
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2619 U$$2756/A1 U$$2663/A2 U$$2756/B1 U$$2663/B2 VGND VGND VPWR VPWR U$$2620/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1907 U$$811/A1 U$$1907/A2 U$$2318/B1 U$$1907/B2 VGND VGND VPWR VPWR U$$1908/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1918 U$$1918/A VGND VGND VPWR VPWR U$$1918/Y sky130_fd_sc_hd__inv_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ _530_/CLK _402_/D VGND VGND VPWR VPWR _402_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1929 U$$1929/A U$$1957/B VGND VGND VPWR VPWR U$$1929/X sky130_fd_sc_hd__xor2_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_333_ _463_/CLK _333_/D VGND VGND VPWR VPWR _333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_264_ _519_/CLK _264_/D VGND VGND VPWR VPWR _264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_195_ _207_/CLK _195_/D VGND VGND VPWR VPWR _195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_95_1 dadda_fa_3_95_1/A dadda_fa_3_95_1/B dadda_fa_3_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_0/CIN dadda_fa_4_95_2/A sky130_fd_sc_hd__fa_1
XFILLER_143_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_72_0 dadda_fa_6_72_0/A dadda_fa_6_72_0/B dadda_fa_6_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_73_0/B dadda_fa_7_72_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_88_0 dadda_fa_3_88_0/A dadda_fa_3_88_0/B dadda_fa_3_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_0/B dadda_fa_4_88_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1025 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater807 U$$2274/B2 VGND VGND VPWR VPWR U$$2262/B2 sky130_fd_sc_hd__buf_4
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4500 U$$938/A1 U$$4388/X U$$4500/B1 U$$4389/X VGND VGND VPWR VPWR U$$4501/A sky130_fd_sc_hd__a22o_1
Xrepeater818 U$$2145/B2 VGND VGND VPWR VPWR U$$2115/B2 sky130_fd_sc_hd__buf_6
XU$$4511 U$$4511/A U$$4511/B VGND VGND VPWR VPWR U$$4511/X sky130_fd_sc_hd__xor2_1
Xrepeater829 U$$2040/B2 VGND VGND VPWR VPWR U$$2052/B2 sky130_fd_sc_hd__buf_6
XFILLER_42_1247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$14 U$$14/A1 U$$8/A2 U$$16/A1 U$$8/B2 VGND VGND VPWR VPWR U$$15/A sky130_fd_sc_hd__a22o_1
XU$$3810 U$$3810/A U$$3836/A VGND VGND VPWR VPWR U$$3810/X sky130_fd_sc_hd__xor2_1
XU$$25 U$$25/A U$$57/B VGND VGND VPWR VPWR U$$25/X sky130_fd_sc_hd__xor2_1
XU$$3821 U$$4506/A1 U$$3703/X U$$4508/A1 U$$3704/X VGND VGND VPWR VPWR U$$3822/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_117_0 U$$3698/Y U$$3832/X U$$3965/X VGND VGND VPWR VPWR dadda_fa_5_118_0/A
+ dadda_fa_5_117_1/A sky130_fd_sc_hd__fa_1
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3832 U$$3832/A U$$3832/B VGND VGND VPWR VPWR U$$3832/X sky130_fd_sc_hd__xor2_1
XU$$36 U$$36/A1 U$$62/A2 U$$38/A1 U$$62/B2 VGND VGND VPWR VPWR U$$37/A sky130_fd_sc_hd__a22o_1
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$47 U$$47/A U$$85/B VGND VGND VPWR VPWR U$$47/X sky130_fd_sc_hd__xor2_1
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3843 U$$3843/A U$$3895/B VGND VGND VPWR VPWR U$$3843/X sky130_fd_sc_hd__xor2_1
XU$$58 U$$58/A1 U$$68/A2 U$$60/A1 U$$68/B2 VGND VGND VPWR VPWR U$$59/A sky130_fd_sc_hd__a22o_1
XU$$3854 U$$4402/A1 U$$3874/A2 U$$4402/B1 U$$3874/B2 VGND VGND VPWR VPWR U$$3855/A
+ sky130_fd_sc_hd__a22o_1
XU$$69 U$$69/A U$$99/B VGND VGND VPWR VPWR U$$69/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_5_4_0 U$$15/X U$$148/X VGND VGND VPWR VPWR dadda_fa_6_5_0/CIN dadda_fa_7_4_0/A
+ sky130_fd_sc_hd__ha_1
XU$$3865 U$$3865/A U$$3949/B VGND VGND VPWR VPWR U$$3865/X sky130_fd_sc_hd__xor2_1
XU$$3876 U$$4287/A1 U$$3910/A2 U$$3876/B1 U$$3910/B2 VGND VGND VPWR VPWR U$$3877/A
+ sky130_fd_sc_hd__a22o_1
XU$$3887 U$$3887/A U$$3917/B VGND VGND VPWR VPWR U$$3887/X sky130_fd_sc_hd__xor2_1
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3898 U$$4444/B1 U$$3910/A2 U$$4446/B1 U$$3910/B2 VGND VGND VPWR VPWR U$$3899/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_16 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_27 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_49 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_90_0 U$$3246/X U$$3379/X U$$3512/X VGND VGND VPWR VPWR dadda_fa_3_91_0/B
+ dadda_fa_3_90_2/B sky130_fd_sc_hd__fa_1
XFILLER_138_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_46_6 U$$2493/X U$$2626/X VGND VGND VPWR VPWR dadda_fa_2_47_3/CIN dadda_fa_3_46_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_87_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_52_5 U$$2372/X U$$2505/X U$$2638/X VGND VGND VPWR VPWR dadda_fa_2_53_2/A
+ dadda_fa_2_52_5/A sky130_fd_sc_hd__fa_1
XFILLER_210_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_45_4 U$$1693/X U$$1826/X U$$1959/X VGND VGND VPWR VPWR dadda_fa_2_46_3/B
+ dadda_fa_2_45_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_15_2 input163/X dadda_fa_4_15_2/B dadda_ha_3_15_0/SUM VGND VGND VPWR VPWR
+ dadda_fa_5_16_0/CIN dadda_fa_5_15_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_184_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1039 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_194 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3106 U$$4476/A1 U$$3110/A2 U$$4478/A1 U$$3110/B2 VGND VGND VPWR VPWR U$$3107/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_1083 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3117 U$$3117/A U$$3121/B VGND VGND VPWR VPWR U$$3117/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3128 _605_/Q U$$3132/A2 _606_/Q U$$3132/B2 VGND VGND VPWR VPWR U$$3129/A sky130_fd_sc_hd__a22o_1
XFILLER_207_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3139 U$$3139/A U$$3145/B VGND VGND VPWR VPWR U$$3139/X sky130_fd_sc_hd__xor2_1
XFILLER_28_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2405 U$$3638/A1 U$$2437/A2 U$$3503/A1 U$$2437/B2 VGND VGND VPWR VPWR U$$2406/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2416 U$$2416/A U$$2436/B VGND VGND VPWR VPWR U$$2416/X sky130_fd_sc_hd__xor2_1
XU$$2427 U$$98/A1 U$$2435/A2 U$$98/B1 U$$2435/B2 VGND VGND VPWR VPWR U$$2428/A sky130_fd_sc_hd__a22o_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2438 U$$2438/A U$$2442/B VGND VGND VPWR VPWR U$$2438/X sky130_fd_sc_hd__xor2_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1704 U$$3485/A1 U$$1710/A2 U$$1843/A1 U$$1710/B2 VGND VGND VPWR VPWR U$$1705/A
+ sky130_fd_sc_hd__a22o_1
XU$$2449 U$$3132/B1 U$$2463/A2 _609_/Q U$$2463/B2 VGND VGND VPWR VPWR U$$2450/A sky130_fd_sc_hd__a22o_1
XU$$1715 U$$1715/A U$$1763/B VGND VGND VPWR VPWR U$$1715/X sky130_fd_sc_hd__xor2_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1726 U$$493/A1 U$$1736/A2 U$$358/A1 U$$1736/B2 VGND VGND VPWR VPWR U$$1727/A sky130_fd_sc_hd__a22o_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1737 U$$1737/A U$$1737/B VGND VGND VPWR VPWR U$$1737/X sky130_fd_sc_hd__xor2_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1748 U$$2431/B1 U$$1768/A2 U$$2435/A1 U$$1768/B2 VGND VGND VPWR VPWR U$$1749/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1759 U$$1759/A U$$1763/B VGND VGND VPWR VPWR U$$1759/X sky130_fd_sc_hd__xor2_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_316_ _445_/CLK _316_/D VGND VGND VPWR VPWR _316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_247_ _504_/CLK _247_/D VGND VGND VPWR VPWR _247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput14 a[21] VGND VGND VPWR VPWR _637_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput25 a[31] VGND VGND VPWR VPWR _647_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_183_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_103_clk _616_/CLK VGND VGND VPWR VPWR _491_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput36 a[41] VGND VGND VPWR VPWR _657_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput47 a[51] VGND VGND VPWR VPWR _667_/D sky130_fd_sc_hd__clkbuf_1
Xinput58 a[61] VGND VGND VPWR VPWR _677_/D sky130_fd_sc_hd__clkbuf_1
X_178_ _189_/CLK _178_/D VGND VGND VPWR VPWR _178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput69 b[13] VGND VGND VPWR VPWR _565_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_526 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_62_4 dadda_fa_2_62_4/A dadda_fa_2_62_4/B dadda_fa_2_62_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/CIN dadda_fa_3_62_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater604 U$$1635/A2 VGND VGND VPWR VPWR U$$1627/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater615 U$$141/X VGND VGND VPWR VPWR U$$263/A2 sky130_fd_sc_hd__buf_4
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater626 U$$1291/A2 VGND VGND VPWR VPWR U$$1295/A2 sky130_fd_sc_hd__buf_4
XFILLER_81_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_55_3 dadda_fa_2_55_3/A dadda_fa_2_55_3/B dadda_fa_2_55_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/B dadda_fa_3_55_3/B sky130_fd_sc_hd__fa_1
XFILLER_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater637 U$$1230/A2 VGND VGND VPWR VPWR U$$1224/A2 sky130_fd_sc_hd__clkbuf_8
XU$$4330 U$$4330/A U$$4334/B VGND VGND VPWR VPWR U$$4330/X sky130_fd_sc_hd__xor2_1
Xrepeater648 U$$928/B2 VGND VGND VPWR VPWR U$$860/B2 sky130_fd_sc_hd__buf_4
Xrepeater659 U$$809/B2 VGND VGND VPWR VPWR U$$819/B2 sky130_fd_sc_hd__buf_8
XU$$4341 U$$4478/A1 U$$4347/A2 U$$4480/A1 U$$4347/B2 VGND VGND VPWR VPWR U$$4342/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4352 U$$4352/A U$$4382/B VGND VGND VPWR VPWR U$$4352/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_48_2 dadda_fa_2_48_2/A dadda_fa_2_48_2/B dadda_fa_2_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/A dadda_fa_3_48_3/A sky130_fd_sc_hd__fa_1
XU$$4363 U$$938/A1 U$$4369/A2 U$$4500/B1 U$$4369/B2 VGND VGND VPWR VPWR U$$4364/A
+ sky130_fd_sc_hd__a22o_1
XU$$4374 U$$4374/A U$$4383/A VGND VGND VPWR VPWR U$$4374/X sky130_fd_sc_hd__xor2_1
XFILLER_77_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4385 U$$4385/A VGND VGND VPWR VPWR U$$4387/B sky130_fd_sc_hd__inv_1
XFILLER_92_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3640 U$$4462/A1 U$$3674/A2 U$$4464/A1 U$$3674/B2 VGND VGND VPWR VPWR U$$3641/A
+ sky130_fd_sc_hd__a22o_1
XU$$3651 U$$3651/A U$$3663/B VGND VGND VPWR VPWR U$$3651/X sky130_fd_sc_hd__xor2_1
XU$$4396 U$$4396/A1 U$$4388/X _555_/Q U$$4438/B2 VGND VGND VPWR VPWR U$$4397/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_25_1 dadda_fa_5_25_1/A dadda_fa_5_25_1/B dadda_fa_5_25_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_26_0/B dadda_fa_7_25_0/A sky130_fd_sc_hd__fa_2
XFILLER_80_502 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3662 _598_/Q U$$3662/A2 U$$3799/B1 U$$3662/B2 VGND VGND VPWR VPWR U$$3663/A sky130_fd_sc_hd__a22o_1
XU$$3673 U$$3673/A _669_/Q VGND VGND VPWR VPWR U$$3673/X sky130_fd_sc_hd__xor2_1
XFILLER_206_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_18_0 dadda_fa_5_18_0/A dadda_fa_5_18_0/B dadda_fa_5_18_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_19_0/A dadda_fa_6_18_0/CIN sky130_fd_sc_hd__fa_2
XU$$3684 U$$4506/A1 U$$3688/A2 U$$4508/A1 U$$3688/B2 VGND VGND VPWR VPWR U$$3685/A
+ sky130_fd_sc_hd__a22o_1
XU$$2950 U$$2950/A U$$2988/B VGND VGND VPWR VPWR U$$2950/X sky130_fd_sc_hd__xor2_1
XU$$3695 U$$3695/A U$$3698/A VGND VGND VPWR VPWR U$$3695/X sky130_fd_sc_hd__xor2_1
XU$$2961 U$$3783/A1 U$$2981/A2 U$$3783/B1 U$$2981/B2 VGND VGND VPWR VPWR U$$2962/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2972 U$$2972/A U$$2972/B VGND VGND VPWR VPWR U$$2972/X sky130_fd_sc_hd__xor2_1
XU$$2983 U$$3805/A1 U$$3005/A2 U$$2983/B1 U$$3005/B2 VGND VGND VPWR VPWR U$$2984/A
+ sky130_fd_sc_hd__a22o_1
XU$$2994 U$$2994/A U$$3000/B VGND VGND VPWR VPWR U$$2994/X sky130_fd_sc_hd__xor2_1
XFILLER_60_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_50_2 U$$905/X U$$1038/X U$$1171/X VGND VGND VPWR VPWR dadda_fa_2_51_1/A
+ dadda_fa_2_50_4/A sky130_fd_sc_hd__fa_1
XFILLER_21_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$806 U$$806/A _627_/Q VGND VGND VPWR VPWR U$$806/X sky130_fd_sc_hd__xor2_1
XU$$817 U$$817/A1 U$$819/A2 U$$817/B1 U$$819/B2 VGND VGND VPWR VPWR U$$818/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_43_1 U$$492/X U$$625/X U$$758/X VGND VGND VPWR VPWR dadda_fa_2_44_3/A
+ dadda_fa_2_43_5/A sky130_fd_sc_hd__fa_1
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$828 U$$828/A1 U$$860/A2 U$$828/B1 U$$860/B2 VGND VGND VPWR VPWR U$$829/A sky130_fd_sc_hd__a22o_1
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$839 U$$839/A U$$859/B VGND VGND VPWR VPWR U$$839/X sky130_fd_sc_hd__xor2_1
XFILLER_73_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_20_0 U$$1429/B input169/X dadda_fa_4_20_0/CIN VGND VGND VPWR VPWR dadda_fa_5_21_0/A
+ dadda_fa_5_20_1/A sky130_fd_sc_hd__fa_1
XFILLER_113_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_36_0 U$$79/X U$$212/X U$$345/X VGND VGND VPWR VPWR dadda_fa_2_37_5/A dadda_fa_2_36_5/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_43_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1706 U$$3157/B1 VGND VGND VPWR VPWR U$$2746/B1 sky130_fd_sc_hd__buf_6
XU$$4491_1824 VGND VGND VPWR VPWR U$$4491_1824/HI U$$4491/B sky130_fd_sc_hd__conb_1
XFILLER_4_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_72_3 dadda_fa_3_72_3/A dadda_fa_3_72_3/B dadda_fa_3_72_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_1/B dadda_fa_4_72_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_65_2 dadda_fa_3_65_2/A dadda_fa_3_65_2/B dadda_fa_3_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_1/A dadda_fa_4_65_2/B sky130_fd_sc_hd__fa_1
XFILLER_117_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_58_1 dadda_fa_3_58_1/A dadda_fa_3_58_1/B dadda_fa_3_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_0/CIN dadda_fa_4_58_2/A sky130_fd_sc_hd__fa_1
XFILLER_117_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_35_0 dadda_fa_6_35_0/A dadda_fa_6_35_0/B dadda_fa_6_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_36_0/B dadda_fa_7_35_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_207_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2202 U$$2611/B1 U$$2242/A2 U$$2478/A1 U$$2242/B2 VGND VGND VPWR VPWR U$$2203/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2213 U$$2213/A U$$2243/B VGND VGND VPWR VPWR U$$2213/X sky130_fd_sc_hd__xor2_1
XU$$2224 U$$3320/A1 U$$2262/A2 U$$3320/B1 U$$2262/B2 VGND VGND VPWR VPWR U$$2225/A
+ sky130_fd_sc_hd__a22o_1
XU$$2235 U$$2235/A U$$2243/B VGND VGND VPWR VPWR U$$2235/X sky130_fd_sc_hd__xor2_1
XU$$2246 U$$4027/A1 U$$2298/A2 _576_/Q U$$2298/B2 VGND VGND VPWR VPWR U$$2247/A sky130_fd_sc_hd__a22o_1
XU$$1501 U$$1501/A U$$1501/B VGND VGND VPWR VPWR U$$1501/X sky130_fd_sc_hd__xor2_1
XU$$1512 U$$1510/B U$$1507/A _638_/Q U$$1507/Y VGND VGND VPWR VPWR U$$1512/X sky130_fd_sc_hd__a22o_2
XFILLER_62_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_952 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2257 U$$2257/A U$$2269/B VGND VGND VPWR VPWR U$$2257/X sky130_fd_sc_hd__xor2_1
XU$$1523 U$$838/A1 U$$1553/A2 U$$840/A1 U$$1553/B2 VGND VGND VPWR VPWR U$$1524/A sky130_fd_sc_hd__a22o_1
XU$$2268 U$$3638/A1 U$$2274/A2 U$$3503/A1 U$$2274/B2 VGND VGND VPWR VPWR U$$2269/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1534 U$$1534/A U$$1562/B VGND VGND VPWR VPWR U$$1534/X sky130_fd_sc_hd__xor2_1
XU$$2279 U$$2279/A U$$2299/B VGND VGND VPWR VPWR U$$2279/X sky130_fd_sc_hd__xor2_1
XU$$1545 U$$449/A1 U$$1561/A2 U$$449/B1 U$$1561/B2 VGND VGND VPWR VPWR U$$1546/A sky130_fd_sc_hd__a22o_1
XU$$1556 U$$1556/A U$$1598/B VGND VGND VPWR VPWR U$$1556/X sky130_fd_sc_hd__xor2_1
XFILLER_187_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1567 U$$745/A1 U$$1587/A2 U$$1843/A1 U$$1587/B2 VGND VGND VPWR VPWR U$$1568/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1578 U$$1578/A U$$1578/B VGND VGND VPWR VPWR U$$1578/X sky130_fd_sc_hd__xor2_1
XFILLER_176_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1589 U$$493/A1 U$$1597/A2 U$$84/A1 U$$1597/B2 VGND VGND VPWR VPWR U$$1590/A sky130_fd_sc_hd__a22o_1
XFILLER_179_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_108_0 dadda_fa_7_108_0/A dadda_fa_7_108_0/B dadda_fa_7_108_0/CIN VGND
+ VGND VPWR VPWR _533_/D _404_/D sky130_fd_sc_hd__fa_1
XFILLER_204_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_112_0_1868 VGND VGND VPWR VPWR dadda_fa_3_112_0/A dadda_fa_3_112_0_1868/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_103_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_60_1 dadda_fa_2_60_1/A dadda_fa_2_60_1/B dadda_fa_2_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_0/CIN dadda_fa_3_60_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater401 U$$765/A2 VGND VGND VPWR VPWR U$$747/A2 sky130_fd_sc_hd__buf_4
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$208 final_adder.U$$703/A final_adder.U$$702/A VGND VGND VPWR VPWR
+ final_adder.U$$296/B sky130_fd_sc_hd__and2_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater412 U$$622/A2 VGND VGND VPWR VPWR U$$632/A2 sky130_fd_sc_hd__buf_8
XFILLER_100_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater423 U$$4251/X VGND VGND VPWR VPWR U$$4335/A2 sky130_fd_sc_hd__buf_6
XFILLER_111_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$219 final_adder.U$$713/A final_adder.U$$585/B1 final_adder.U$$219/B1
+ VGND VGND VPWR VPWR final_adder.U$$219/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_2_53_0 dadda_fa_2_53_0/A dadda_fa_2_53_0/B dadda_fa_2_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_0/B dadda_fa_3_53_2/B sky130_fd_sc_hd__fa_2
XFILLER_38_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater434 U$$4114/X VGND VGND VPWR VPWR U$$4244/A2 sky130_fd_sc_hd__buf_4
XFILLER_211_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater445 U$$4/X VGND VGND VPWR VPWR U$$98/A2 sky130_fd_sc_hd__buf_4
Xrepeater456 U$$3840/X VGND VGND VPWR VPWR U$$3932/A2 sky130_fd_sc_hd__buf_4
Xrepeater467 U$$3805/A2 VGND VGND VPWR VPWR U$$3777/A2 sky130_fd_sc_hd__buf_6
Xrepeater478 U$$3497/A2 VGND VGND VPWR VPWR U$$3479/A2 sky130_fd_sc_hd__buf_8
XU$$4160 U$$4160/A1 U$$4174/A2 U$$4160/B1 U$$4174/B2 VGND VGND VPWR VPWR U$$4161/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater489 U$$3378/A2 VGND VGND VPWR VPWR U$$3356/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_66_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4171 U$$4171/A U$$4215/B VGND VGND VPWR VPWR U$$4171/X sky130_fd_sc_hd__xor2_1
XU$$4182 U$$4317/B1 U$$4182/A2 U$$4184/A1 U$$4182/B2 VGND VGND VPWR VPWR U$$4183/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4193 U$$4193/A U$$4197/B VGND VGND VPWR VPWR U$$4193/X sky130_fd_sc_hd__xor2_1
XFILLER_129_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3470 U$$3470/A U$$3506/B VGND VGND VPWR VPWR U$$3470/X sky130_fd_sc_hd__xor2_1
XFILLER_92_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3481 U$$3618/A1 U$$3519/A2 _577_/Q U$$3519/B2 VGND VGND VPWR VPWR U$$3482/A sky130_fd_sc_hd__a22o_1
XU$$3492 U$$3492/A U$$3520/B VGND VGND VPWR VPWR U$$3492/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_7_0 U$$21/X U$$154/X U$$287/X VGND VGND VPWR VPWR dadda_fa_6_8_0/A dadda_fa_6_7_0/CIN
+ sky130_fd_sc_hd__fa_2
XFILLER_94_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2780 U$$451/A1 U$$2812/A2 U$$3876/B1 U$$2812/B2 VGND VGND VPWR VPWR U$$2781/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2791 U$$2791/A U$$2795/B VGND VGND VPWR VPWR U$$2791/X sky130_fd_sc_hd__xor2_1
XFILLER_179_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_1084 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_418 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_82_2 dadda_fa_4_82_2/A dadda_fa_4_82_2/B dadda_fa_4_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/CIN dadda_fa_5_82_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_75_1 dadda_fa_4_75_1/A dadda_fa_4_75_1/B dadda_fa_4_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/B dadda_fa_5_75_1/B sky130_fd_sc_hd__fa_1
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_52_0 dadda_fa_7_52_0/A dadda_fa_7_52_0/B dadda_fa_7_52_0/CIN VGND VGND
+ VPWR VPWR _477_/D _348_/D sky130_fd_sc_hd__fa_1
XFILLER_0_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_68_0 dadda_fa_4_68_0/A dadda_fa_4_68_0/B dadda_fa_4_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/A dadda_fa_5_68_1/A sky130_fd_sc_hd__fa_1
XFILLER_88_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput204 c[52] VGND VGND VPWR VPWR input204/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput215 c[62] VGND VGND VPWR VPWR input215/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput226 c[72] VGND VGND VPWR VPWR input226/X sky130_fd_sc_hd__buf_2
XTAP_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 c[82] VGND VGND VPWR VPWR input237/X sky130_fd_sc_hd__buf_2
XTAP_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput248 c[92] VGND VGND VPWR VPWR input248/X sky130_fd_sc_hd__clkbuf_4
XTAP_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$720 final_adder.U$$720/A final_adder.U$$720/B VGND VGND VPWR VPWR
+ _266_/D sky130_fd_sc_hd__xor2_1
XTAP_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$731 final_adder.U$$731/A final_adder.U$$731/B VGND VGND VPWR VPWR
+ _277_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$742 final_adder.U$$742/A final_adder.U$$742/B VGND VGND VPWR VPWR
+ _288_/D sky130_fd_sc_hd__xor2_4
X_650_ _660_/CLK _650_/D VGND VGND VPWR VPWR _650_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$603 U$$603/A U$$613/B VGND VGND VPWR VPWR U$$603/X sky130_fd_sc_hd__xor2_1
XFILLER_5_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$614 U$$614/A1 U$$616/A2 U$$614/B1 U$$616/B2 VGND VGND VPWR VPWR U$$615/A sky130_fd_sc_hd__a22o_1
Xrepeater990 U$$3121/B VGND VGND VPWR VPWR U$$3133/B sky130_fd_sc_hd__buf_6
XU$$625 U$$625/A U$$669/B VGND VGND VPWR VPWR U$$625/X sky130_fd_sc_hd__xor2_1
X_581_ _582_/CLK _581_/D VGND VGND VPWR VPWR _581_/Q sky130_fd_sc_hd__dfxtp_1
XU$$636 U$$910/A1 U$$650/A2 U$$912/A1 U$$650/B2 VGND VGND VPWR VPWR U$$637/A sky130_fd_sc_hd__a22o_1
XFILLER_29_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$647 U$$647/A U$$651/B VGND VGND VPWR VPWR U$$647/X sky130_fd_sc_hd__xor2_1
XFILLER_205_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$658 U$$658/A1 U$$682/A2 U$$658/B1 U$$682/B2 VGND VGND VPWR VPWR U$$659/A sky130_fd_sc_hd__a22o_1
XU$$669 U$$669/A U$$669/B VGND VGND VPWR VPWR U$$669/X sky130_fd_sc_hd__xor2_1
XFILLER_189_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1503 U$$467/B1 VGND VGND VPWR VPWR U$$2796/B1 sky130_fd_sc_hd__buf_4
Xrepeater1514 U$$4440/A1 VGND VGND VPWR VPWR U$$4027/B1 sky130_fd_sc_hd__buf_8
Xrepeater1525 U$$4160/B1 VGND VGND VPWR VPWR U$$3751/A1 sky130_fd_sc_hd__buf_4
Xrepeater1536 U$$3475/A1 VGND VGND VPWR VPWR U$$733/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_180_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1547 _572_/Q VGND VGND VPWR VPWR U$$4156/B1 sky130_fd_sc_hd__buf_6
XFILLER_99_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1558 U$$3056/B1 VGND VGND VPWR VPWR U$$866/A1 sky130_fd_sc_hd__buf_8
Xrepeater1569 _569_/Q VGND VGND VPWR VPWR U$$4426/A1 sky130_fd_sc_hd__buf_6
XFILLER_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_70_0 dadda_fa_3_70_0/A dadda_fa_3_70_0/B dadda_fa_3_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_0/B dadda_fa_4_70_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2010 U$$229/A1 U$$2010/A2 U$$2832/B1 U$$2010/B2 VGND VGND VPWR VPWR U$$2011/A
+ sky130_fd_sc_hd__a22o_1
XU$$2021 U$$2021/A U$$2029/B VGND VGND VPWR VPWR U$$2021/X sky130_fd_sc_hd__xor2_1
XFILLER_130_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2032 U$$2717/A1 U$$2038/A2 U$$2171/A1 U$$2038/B2 VGND VGND VPWR VPWR U$$2033/A
+ sky130_fd_sc_hd__a22o_1
XU$$2043 U$$2043/A U$$2043/B VGND VGND VPWR VPWR U$$2043/X sky130_fd_sc_hd__xor2_1
XU$$2054 U$$2054/A VGND VGND VPWR VPWR U$$2054/Y sky130_fd_sc_hd__inv_1
XFILLER_62_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1320 U$$1320/A U$$1356/B VGND VGND VPWR VPWR U$$1320/X sky130_fd_sc_hd__xor2_1
XU$$2065 U$$2611/B1 U$$2115/A2 U$$2478/A1 U$$2115/B2 VGND VGND VPWR VPWR U$$2066/A
+ sky130_fd_sc_hd__a22o_1
XU$$1331 U$$2838/A1 U$$1237/X U$$2838/B1 U$$1238/X VGND VGND VPWR VPWR U$$1332/A sky130_fd_sc_hd__a22o_1
XU$$2076 U$$2076/A U$$2108/B VGND VGND VPWR VPWR U$$2076/X sky130_fd_sc_hd__xor2_1
XU$$2087 U$$32/A1 U$$2129/A2 U$$993/A1 U$$2129/B2 VGND VGND VPWR VPWR U$$2088/A sky130_fd_sc_hd__a22o_1
XU$$1342 U$$1342/A U$$1369/A VGND VGND VPWR VPWR U$$1342/X sky130_fd_sc_hd__xor2_1
XU$$1353 U$$2721/B1 U$$1355/A2 U$$2725/A1 U$$1355/B2 VGND VGND VPWR VPWR U$$1354/A
+ sky130_fd_sc_hd__a22o_1
XU$$2098 U$$2098/A U$$2110/B VGND VGND VPWR VPWR U$$2098/X sky130_fd_sc_hd__xor2_1
XU$$1364 U$$1364/A U$$1368/B VGND VGND VPWR VPWR U$$1364/X sky130_fd_sc_hd__xor2_1
XFILLER_95_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1375 U$$1373/B _635_/Q _636_/Q U$$1370/Y VGND VGND VPWR VPWR U$$1375/X sky130_fd_sc_hd__a22o_4
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1386 U$$973/B1 U$$1424/A2 U$$2756/B1 U$$1424/B2 VGND VGND VPWR VPWR U$$1387/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1397 U$$1397/A U$$1425/B VGND VGND VPWR VPWR U$$1397/X sky130_fd_sc_hd__xor2_1
XFILLER_149_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_92_1 dadda_fa_5_92_1/A dadda_fa_5_92_1/B dadda_fa_5_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_93_0/B dadda_fa_7_92_0/A sky130_fd_sc_hd__fa_1
XFILLER_157_982 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_85_0 dadda_fa_5_85_0/A dadda_fa_5_85_0/B dadda_fa_5_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_86_0/A dadda_fa_6_85_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_190_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_77_7 U$$4151/X U$$4284/X U$$4417/X VGND VGND VPWR VPWR dadda_fa_2_78_2/CIN
+ dadda_fa_2_77_5/CIN sky130_fd_sc_hd__fa_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_309 _236_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_92_clk _628_/CLK VGND VGND VPWR VPWR _642_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$60 _484_/Q _356_/Q VGND VGND VPWR VPWR final_adder.U$$555/B1 final_adder.U$$682/A
+ sky130_fd_sc_hd__ha_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$71 _495_/Q _367_/Q VGND VGND VPWR VPWR final_adder.U$$199/B1 final_adder.U$$693/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$82 _506_/Q _378_/Q VGND VGND VPWR VPWR final_adder.U$$577/B1 final_adder.U$$704/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$93 _517_/Q _389_/Q VGND VGND VPWR VPWR final_adder.U$$221/B1 final_adder.U$$715/A
+ sky130_fd_sc_hd__ha_1
XFILLER_41_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_101_2 dadda_fa_3_101_2/A dadda_fa_3_101_2/B dadda_fa_3_101_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_102_1/A dadda_fa_4_101_2/B sky130_fd_sc_hd__fa_1
XFILLER_150_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_495 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_65_5 U$$2132/X U$$2265/X U$$2398/X VGND VGND VPWR VPWR dadda_fa_1_66_7/A
+ dadda_fa_2_65_0/A sky130_fd_sc_hd__fa_1
XTAP_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_115_0 dadda_fa_6_115_0/A dadda_fa_6_115_0/B dadda_fa_6_115_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_116_0/B dadda_fa_7_115_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$400 U$$674/A1 U$$408/A2 U$$676/A1 U$$408/B2 VGND VGND VPWR VPWR U$$401/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$561 final_adder.U$$688/A final_adder.U$$688/B final_adder.U$$561/B1
+ VGND VGND VPWR VPWR final_adder.U$$689/B sky130_fd_sc_hd__a21o_1
XTAP_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_633_ _633_/CLK _633_/D VGND VGND VPWR VPWR _633_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$411 U$$411/A VGND VGND VPWR VPWR U$$411/Y sky130_fd_sc_hd__inv_1
XTAP_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_35_3 dadda_fa_3_35_3/A dadda_fa_3_35_3/B dadda_fa_3_35_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_1/B dadda_fa_4_35_2/CIN sky130_fd_sc_hd__fa_1
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$422 U$$422/A U$$452/B VGND VGND VPWR VPWR U$$422/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$583 final_adder.U$$710/A final_adder.U$$710/B final_adder.U$$583/B1
+ VGND VGND VPWR VPWR final_adder.U$$711/B sky130_fd_sc_hd__a21o_1
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$433 U$$707/A1 U$$457/A2 U$$22/B1 U$$457/B2 VGND VGND VPWR VPWR U$$434/A sky130_fd_sc_hd__a22o_1
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_clk _628_/CLK VGND VGND VPWR VPWR _550_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$444 U$$444/A U$$452/B VGND VGND VPWR VPWR U$$444/X sky130_fd_sc_hd__xor2_1
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$455 U$$42/B1 U$$457/A2 U$$729/B1 U$$457/B2 VGND VGND VPWR VPWR U$$456/A sky130_fd_sc_hd__a22o_1
XFILLER_72_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_564_ _569_/CLK _564_/D VGND VGND VPWR VPWR _564_/Q sky130_fd_sc_hd__dfxtp_4
Xdadda_fa_3_28_2 dadda_fa_3_28_2/A dadda_fa_3_28_2/B dadda_fa_3_28_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_29_1/A dadda_fa_4_28_2/B sky130_fd_sc_hd__fa_1
XFILLER_189_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$466 U$$466/A U$$500/B VGND VGND VPWR VPWR U$$466/X sky130_fd_sc_hd__xor2_1
XU$$477 U$$614/A1 U$$483/A2 U$$614/B1 U$$483/B2 VGND VGND VPWR VPWR U$$478/A sky130_fd_sc_hd__a22o_1
XFILLER_44_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$488 U$$488/A U$$532/B VGND VGND VPWR VPWR U$$488/X sky130_fd_sc_hd__xor2_1
XFILLER_32_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$499 U$$634/B1 U$$499/A2 U$$501/A1 U$$499/B2 VGND VGND VPWR VPWR U$$500/A sky130_fd_sc_hd__a22o_1
XFILLER_38_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_495_ _495_/CLK _495_/D VGND VGND VPWR VPWR _495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_396 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_610 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1300 U$$2983/B1 VGND VGND VPWR VPWR U$$791/B1 sky130_fd_sc_hd__buf_6
XFILLER_172_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1311 U$$3942/A1 VGND VGND VPWR VPWR U$$4353/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1322 _600_/Q VGND VGND VPWR VPWR U$$3529/A1 sky130_fd_sc_hd__buf_6
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1333 _598_/Q VGND VGND VPWR VPWR U$$3386/B1 sky130_fd_sc_hd__buf_4
XFILLER_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1344 U$$4206/B1 VGND VGND VPWR VPWR U$$4482/A1 sky130_fd_sc_hd__buf_4
Xrepeater1355 U$$916/A1 VGND VGND VPWR VPWR U$$914/B1 sky130_fd_sc_hd__buf_4
XFILLER_125_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1366 _594_/Q VGND VGND VPWR VPWR U$$3380/A1 sky130_fd_sc_hd__buf_6
XFILLER_4_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1377 U$$4198/B1 VGND VGND VPWR VPWR U$$4472/B1 sky130_fd_sc_hd__buf_6
Xrepeater1388 U$$2415/A1 VGND VGND VPWR VPWR U$$84/B1 sky130_fd_sc_hd__buf_6
Xrepeater1399 U$$3372/A1 VGND VGND VPWR VPWR U$$358/A1 sky130_fd_sc_hd__buf_4
XFILLER_171_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_2_31_4 U$$1665/X U$$1798/X VGND VGND VPWR VPWR dadda_fa_3_32_2/A dadda_fa_4_31_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_94_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_755 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_7_1_0 U$$9/X input168/X VGND VGND VPWR VPWR _426_/D _297_/D sky130_fd_sc_hd__ha_1
XFILLER_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_671 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_74_clk _634_/CLK VGND VGND VPWR VPWR _515_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_2_30_2 U$$865/X U$$998/X U$$1131/X VGND VGND VPWR VPWR dadda_fa_3_31_1/CIN
+ dadda_fa_3_30_3/B sky130_fd_sc_hd__fa_1
XFILLER_211_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_814 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1150 U$$463/B1 U$$1150/A2 U$$330/A1 U$$1150/B2 VGND VGND VPWR VPWR U$$1151/A sky130_fd_sc_hd__a22o_1
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1161 U$$1161/A U$$1191/B VGND VGND VPWR VPWR U$$1161/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1172 U$$898/A1 U$$1176/A2 U$$78/A1 U$$1176/B2 VGND VGND VPWR VPWR U$$1173/A sky130_fd_sc_hd__a22o_1
XFILLER_204_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1183 U$$1183/A U$$1225/B VGND VGND VPWR VPWR U$$1183/X sky130_fd_sc_hd__xor2_1
XU$$1194 U$$2838/A1 U$$1194/A2 U$$2838/B1 U$$1194/B2 VGND VGND VPWR VPWR U$$1195/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_82_5 U$$3230/X U$$3363/X U$$3496/X VGND VGND VPWR VPWR dadda_fa_2_83_3/A
+ dadda_fa_2_82_5/B sky130_fd_sc_hd__fa_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_75_4 U$$3216/X U$$3349/X U$$3482/X VGND VGND VPWR VPWR dadda_fa_2_76_1/CIN
+ dadda_fa_2_75_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_3 U$$3734/X U$$3867/X U$$4000/X VGND VGND VPWR VPWR dadda_fa_2_69_1/B
+ dadda_fa_2_68_4/B sky130_fd_sc_hd__fa_1
XFILLER_105_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_45_2 dadda_fa_4_45_2/A dadda_fa_4_45_2/B dadda_fa_4_45_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/CIN dadda_fa_5_45_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_85_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_1 dadda_fa_4_38_1/A dadda_fa_4_38_1/B dadda_fa_4_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/B dadda_fa_5_38_1/B sky130_fd_sc_hd__fa_1
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_106 _287_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_7_15_0 dadda_fa_7_15_0/A dadda_fa_7_15_0/B dadda_fa_7_15_0/CIN VGND VGND
+ VPWR VPWR _440_/D _311_/D sky130_fd_sc_hd__fa_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_65_clk _535_/CLK VGND VGND VPWR VPWR _530_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_117 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_199_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_128 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_139 _290_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_26 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_280_ _523_/CLK _280_/D VGND VGND VPWR VPWR _280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_70_3 U$$1610/X U$$1743/X U$$1876/X VGND VGND VPWR VPWR dadda_fa_1_71_7/B
+ dadda_fa_1_70_8/CIN sky130_fd_sc_hd__fa_1
XTAP_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_2 U$$931/X U$$1064/X U$$1197/X VGND VGND VPWR VPWR dadda_fa_1_64_6/A
+ dadda_fa_1_63_8/A sky130_fd_sc_hd__fa_1
XTAP_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_917 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_40_1 dadda_fa_3_40_1/A dadda_fa_3_40_1/B dadda_fa_3_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_0/CIN dadda_fa_4_40_2/A sky130_fd_sc_hd__fa_1
XTAP_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_56_1 U$$518/X U$$651/X U$$784/X VGND VGND VPWR VPWR dadda_fa_1_57_7/CIN
+ dadda_fa_1_56_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_56_clk _535_/CLK VGND VGND VPWR VPWR _613_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_33_0 input183/X dadda_fa_3_33_0/B dadda_fa_3_33_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_34_0/B dadda_fa_4_33_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$230 U$$230/A U$$232/B VGND VGND VPWR VPWR U$$230/X sky130_fd_sc_hd__xor2_1
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_616_ _616_/CLK _616_/D VGND VGND VPWR VPWR U$$1/A sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$391 final_adder.U$$354/B final_adder.U$$638/B final_adder.U$$325/X
+ VGND VGND VPWR VPWR final_adder.U$$646/B sky130_fd_sc_hd__a21o_2
XFILLER_205_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$241 U$$650/B1 U$$249/A2 U$$515/B1 U$$249/B2 VGND VGND VPWR VPWR U$$242/A sky130_fd_sc_hd__a22o_1
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$252 U$$252/A U$$264/B VGND VGND VPWR VPWR U$$252/X sky130_fd_sc_hd__xor2_1
XFILLER_205_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$263 U$$674/A1 U$$263/A2 U$$676/A1 U$$263/B2 VGND VGND VPWR VPWR U$$264/A sky130_fd_sc_hd__a22o_1
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_899 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$274 _619_/Q VGND VGND VPWR VPWR U$$274/Y sky130_fd_sc_hd__inv_1
XFILLER_45_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$285 U$$285/A U$$319/B VGND VGND VPWR VPWR U$$285/X sky130_fd_sc_hd__xor2_1
X_547_ _547_/CLK _547_/D VGND VGND VPWR VPWR _547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$296 U$$707/A1 U$$308/A2 U$$22/B1 U$$308/B2 VGND VGND VPWR VPWR U$$297/A sky130_fd_sc_hd__a22o_1
XFILLER_60_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_478_ _478_/CLK _478_/D VGND VGND VPWR VPWR _478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_1216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2 U$$2/A VGND VGND VPWR VPWR U$$2/Y sky130_fd_sc_hd__inv_1
XFILLER_69_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput305 _196_/Q VGND VGND VPWR VPWR o[28] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_4 input248/X dadda_fa_2_92_4/B dadda_fa_2_92_4/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_93_1/CIN dadda_fa_3_92_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_127_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1130 U$$935/B VGND VGND VPWR VPWR U$$929/B sky130_fd_sc_hd__buf_6
XFILLER_58_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput316 _206_/Q VGND VGND VPWR VPWR o[38] sky130_fd_sc_hd__buf_2
Xoutput327 _216_/Q VGND VGND VPWR VPWR o[48] sky130_fd_sc_hd__buf_2
Xrepeater1141 U$$766/B VGND VGND VPWR VPWR U$$748/B sky130_fd_sc_hd__buf_6
Xoutput338 _226_/Q VGND VGND VPWR VPWR o[58] sky130_fd_sc_hd__buf_2
XFILLER_141_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1152 U$$669/B VGND VGND VPWR VPWR U$$627/B sky130_fd_sc_hd__buf_8
Xoutput349 _236_/Q VGND VGND VPWR VPWR o[68] sky130_fd_sc_hd__buf_2
Xrepeater1163 _623_/Q VGND VGND VPWR VPWR U$$547/A sky130_fd_sc_hd__buf_8
Xdadda_fa_2_85_3 dadda_fa_2_85_3/A dadda_fa_2_85_3/B dadda_fa_2_85_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/B dadda_fa_3_85_3/B sky130_fd_sc_hd__fa_1
Xrepeater1174 U$$226/B VGND VGND VPWR VPWR U$$196/B sky130_fd_sc_hd__buf_6
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1185 U$$85/B VGND VGND VPWR VPWR U$$9/B sky130_fd_sc_hd__buf_4
XFILLER_4_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1196 U$$3285/A1 VGND VGND VPWR VPWR U$$4516/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_206_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_78_2 dadda_fa_2_78_2/A dadda_fa_2_78_2/B dadda_fa_2_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/A dadda_fa_3_78_3/A sky130_fd_sc_hd__fa_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_55_1 dadda_fa_5_55_1/A dadda_fa_5_55_1/B dadda_fa_5_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_56_0/B dadda_fa_7_55_0/A sky130_fd_sc_hd__fa_1
XFILLER_136_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_48_0 dadda_fa_5_48_0/A dadda_fa_5_48_0/B dadda_fa_5_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_49_0/A dadda_fa_6_48_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_ha_2_22_0 U$$51/X U$$184/X VGND VGND VPWR VPWR dadda_fa_3_23_3/CIN dadda_fa_4_22_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_110_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_clk _369_/CLK VGND VGND VPWR VPWR _253_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_674 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_101_1 U$$3002/X U$$3135/X U$$3268/X VGND VGND VPWR VPWR dadda_fa_3_102_2/A
+ dadda_fa_3_101_3/B sky130_fd_sc_hd__fa_1
XFILLER_63_482 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_122_0 U$$4241/X U$$4374/X U$$4507/X VGND VGND VPWR VPWR dadda_fa_6_123_0/A
+ dadda_fa_6_122_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_52_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_80_2 U$$1896/X U$$2029/X U$$2162/X VGND VGND VPWR VPWR dadda_fa_2_81_1/B
+ dadda_fa_2_80_4/A sky130_fd_sc_hd__fa_1
XFILLER_120_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_73_1 U$$2281/X U$$2414/X U$$2547/X VGND VGND VPWR VPWR dadda_fa_2_74_0/CIN
+ dadda_fa_2_73_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_50_0 dadda_fa_4_50_0/A dadda_fa_4_50_0/B dadda_fa_4_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/A dadda_fa_5_50_1/A sky130_fd_sc_hd__fa_1
XFILLER_86_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_66_0 U$$2533/X U$$2666/X U$$2799/X VGND VGND VPWR VPWR dadda_fa_2_67_0/B
+ dadda_fa_2_66_3/B sky130_fd_sc_hd__fa_1
XFILLER_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_clk _479_/CLK VGND VGND VPWR VPWR _484_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2609 U$$2609/A1 U$$2697/A2 U$$2611/A1 U$$2697/B2 VGND VGND VPWR VPWR U$$2610/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1908 U$$1908/A U$$1918/A VGND VGND VPWR VPWR U$$1908/X sky130_fd_sc_hd__xor2_1
XFILLER_148_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1919 _644_/Q VGND VGND VPWR VPWR U$$1921/B sky130_fd_sc_hd__inv_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_401_ _530_/CLK _401_/D VGND VGND VPWR VPWR _401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_332_ _463_/CLK _332_/D VGND VGND VPWR VPWR _332_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_263_ _519_/CLK _263_/D VGND VGND VPWR VPWR _263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_194_ _207_/CLK _194_/D VGND VGND VPWR VPWR _194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4455_1806 VGND VGND VPWR VPWR U$$4455_1806/HI U$$4455/B sky130_fd_sc_hd__conb_1
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_95_2 dadda_fa_3_95_2/A dadda_fa_3_95_2/B dadda_fa_3_95_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_1/A dadda_fa_4_95_2/B sky130_fd_sc_hd__fa_1
XFILLER_136_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_88_1 dadda_fa_3_88_1/A dadda_fa_3_88_1/B dadda_fa_3_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_0/CIN dadda_fa_4_88_2/A sky130_fd_sc_hd__fa_1
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_65_0 dadda_fa_6_65_0/A dadda_fa_6_65_0/B dadda_fa_6_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_66_0/B dadda_fa_7_65_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$6_1841 VGND VGND VPWR VPWR U$$6_1841/HI U$$6/A1 sky130_fd_sc_hd__conb_1
Xrepeater808 U$$2248/B2 VGND VGND VPWR VPWR U$$2242/B2 sky130_fd_sc_hd__clkbuf_4
Xrepeater819 U$$2169/B2 VGND VGND VPWR VPWR U$$2145/B2 sky130_fd_sc_hd__buf_6
XU$$4501 U$$4501/A U$$4501/B VGND VGND VPWR VPWR U$$4501/X sky130_fd_sc_hd__xor2_1
XFILLER_77_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4512 U$$4512/A1 U$$4388/X U$$4514/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4513/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3800 U$$3800/A U$$3800/B VGND VGND VPWR VPWR U$$3800/X sky130_fd_sc_hd__xor2_1
XFILLER_65_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$15 U$$15/A U$$9/B VGND VGND VPWR VPWR U$$15/X sky130_fd_sc_hd__xor2_1
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3811 U$$4222/A1 U$$3823/A2 U$$4087/A1 U$$3823/B2 VGND VGND VPWR VPWR U$$3812/A
+ sky130_fd_sc_hd__a22o_1
XU$$26 U$$26/A1 U$$52/A2 U$$28/A1 U$$52/B2 VGND VGND VPWR VPWR U$$27/A sky130_fd_sc_hd__a22o_1
XFILLER_92_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3822 U$$3822/A U$$3835/A VGND VGND VPWR VPWR U$$3822/X sky130_fd_sc_hd__xor2_1
XU$$37 U$$37/A U$$3/A VGND VGND VPWR VPWR U$$37/X sky130_fd_sc_hd__xor2_1
XU$$4388_1771 VGND VGND VPWR VPWR U$$4388_1771/HI U$$4388/A2 sky130_fd_sc_hd__conb_1
Xdadda_fa_4_117_1 U$$4098/X U$$4231/X U$$4364/X VGND VGND VPWR VPWR dadda_fa_5_118_0/B
+ dadda_fa_5_117_1/B sky130_fd_sc_hd__fa_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_29_clk _432_/CLK VGND VGND VPWR VPWR _478_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3833 U$$4105/B1 U$$3833/A2 U$$3833/B1 U$$3833/B2 VGND VGND VPWR VPWR U$$3834/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$48 U$$48/A1 U$$8/A2 U$$48/B1 U$$8/B2 VGND VGND VPWR VPWR U$$49/A sky130_fd_sc_hd__a22o_1
XU$$3844 U$$3844/A1 U$$3874/A2 _553_/Q U$$3874/B2 VGND VGND VPWR VPWR U$$3845/A sky130_fd_sc_hd__a22o_1
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$59 U$$59/A U$$93/B VGND VGND VPWR VPWR U$$59/X sky130_fd_sc_hd__xor2_1
XFILLER_18_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3855 U$$3855/A U$$3873/B VGND VGND VPWR VPWR U$$3855/X sky130_fd_sc_hd__xor2_1
XFILLER_80_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3866 U$$4003/A1 U$$3958/A2 _564_/Q U$$3958/B2 VGND VGND VPWR VPWR U$$3867/A sky130_fd_sc_hd__a22o_1
XU$$3877 U$$3877/A U$$3933/B VGND VGND VPWR VPWR U$$3877/X sky130_fd_sc_hd__xor2_1
XFILLER_166_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3888 U$$4160/B1 U$$3916/A2 U$$4027/A1 U$$3916/B2 VGND VGND VPWR VPWR U$$3889/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3899 U$$3899/A U$$3933/B VGND VGND VPWR VPWR U$$3899/X sky130_fd_sc_hd__xor2_1
XFILLER_61_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_17 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_28 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _283_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_90_1 U$$3645/X U$$3778/X U$$3911/X VGND VGND VPWR VPWR dadda_fa_3_91_0/CIN
+ dadda_fa_3_90_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_127_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_83_0 U$$4163/X U$$4296/X U$$4429/X VGND VGND VPWR VPWR dadda_fa_3_84_0/B
+ dadda_fa_3_83_2/B sky130_fd_sc_hd__fa_1
XFILLER_142_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_52_6 U$$2771/X U$$2904/X U$$3037/X VGND VGND VPWR VPWR dadda_fa_2_53_2/B
+ dadda_fa_2_52_5/B sky130_fd_sc_hd__fa_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_4_0 dadda_fa_7_4_0/A dadda_fa_7_4_0/B dadda_fa_7_4_0/CIN VGND VGND VPWR
+ VPWR _429_/D _300_/D sky130_fd_sc_hd__fa_1
XFILLER_110_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_82_0 dadda_fa_7_82_0/A dadda_fa_7_82_0/B dadda_fa_7_82_0/CIN VGND VGND
+ VPWR VPWR _507_/D _378_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_98_0 dadda_fa_4_98_0/A dadda_fa_4_98_0/B dadda_fa_4_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/A dadda_fa_5_98_1/A sky130_fd_sc_hd__fa_1
XFILLER_165_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3107 U$$3107/A U$$3107/B VGND VGND VPWR VPWR U$$3107/X sky130_fd_sc_hd__xor2_1
XFILLER_207_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3118 U$$3253/B1 U$$3120/A2 U$$3255/B1 U$$3120/B2 VGND VGND VPWR VPWR U$$3119/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1095 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3129 U$$3129/A U$$3133/B VGND VGND VPWR VPWR U$$3129/X sky130_fd_sc_hd__xor2_1
XFILLER_35_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2406 U$$2406/A U$$2442/B VGND VGND VPWR VPWR U$$2406/X sky130_fd_sc_hd__xor2_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2417 U$$910/A1 U$$2423/A2 U$$912/A1 U$$2423/B2 VGND VGND VPWR VPWR U$$2418/A sky130_fd_sc_hd__a22o_1
XU$$2428 U$$2428/A U$$2436/B VGND VGND VPWR VPWR U$$2428/X sky130_fd_sc_hd__xor2_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2439 U$$4357/A1 U$$2333/X U$$4494/B1 U$$2334/X VGND VGND VPWR VPWR U$$2440/A sky130_fd_sc_hd__a22o_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1705 U$$1705/A U$$1711/B VGND VGND VPWR VPWR U$$1705/X sky130_fd_sc_hd__xor2_1
XFILLER_55_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1716 U$$2947/B1 U$$1718/A2 U$$896/A1 U$$1718/B2 VGND VGND VPWR VPWR U$$1717/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1727 U$$1727/A U$$1737/B VGND VGND VPWR VPWR U$$1727/X sky130_fd_sc_hd__xor2_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1738 U$$2832/B1 U$$1740/A2 U$$3245/B1 U$$1740/B2 VGND VGND VPWR VPWR U$$1739/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1749 U$$1749/A U$$1773/B VGND VGND VPWR VPWR U$$1749/X sky130_fd_sc_hd__xor2_1
XFILLER_202_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_315_ _443_/CLK _315_/D VGND VGND VPWR VPWR _315_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_246_ _504_/CLK _246_/D VGND VGND VPWR VPWR _246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput15 a[22] VGND VGND VPWR VPWR _638_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput26 a[32] VGND VGND VPWR VPWR _648_/D sky130_fd_sc_hd__clkbuf_1
Xinput37 a[42] VGND VGND VPWR VPWR _658_/D sky130_fd_sc_hd__clkbuf_1
Xinput48 a[52] VGND VGND VPWR VPWR _668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput59 a[62] VGND VGND VPWR VPWR _678_/D sky130_fd_sc_hd__clkbuf_1
X_177_ _179_/CLK _177_/D VGND VGND VPWR VPWR _177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_62_5 dadda_fa_2_62_5/A dadda_fa_2_62_5/B dadda_fa_2_62_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_2/A dadda_fa_4_62_0/A sky130_fd_sc_hd__fa_2
Xrepeater605 U$$1635/A2 VGND VGND VPWR VPWR U$$1587/A2 sky130_fd_sc_hd__buf_6
Xrepeater616 U$$1458/A2 VGND VGND VPWR VPWR U$$1424/A2 sky130_fd_sc_hd__buf_4
Xrepeater627 U$$1323/A2 VGND VGND VPWR VPWR U$$1291/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_55_4 dadda_fa_2_55_4/A dadda_fa_2_55_4/B dadda_fa_2_55_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/CIN dadda_fa_3_55_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater638 U$$1208/A2 VGND VGND VPWR VPWR U$$1230/A2 sky130_fd_sc_hd__buf_8
XU$$4320 U$$4320/A U$$4322/B VGND VGND VPWR VPWR U$$4320/X sky130_fd_sc_hd__xor2_1
Xrepeater649 U$$827/X VGND VGND VPWR VPWR U$$928/B2 sky130_fd_sc_hd__buf_4
XU$$4331 U$$4468/A1 U$$4335/A2 U$$4470/A1 U$$4333/B2 VGND VGND VPWR VPWR U$$4332/A
+ sky130_fd_sc_hd__a22o_1
XU$$4342 U$$4342/A U$$4348/B VGND VGND VPWR VPWR U$$4342/X sky130_fd_sc_hd__xor2_1
XFILLER_77_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4353 U$$4353/A1 U$$4369/A2 U$$4490/B1 U$$4369/B2 VGND VGND VPWR VPWR U$$4354/A
+ sky130_fd_sc_hd__a22o_1
XU$$4364 U$$4364/A U$$4384/A VGND VGND VPWR VPWR U$$4364/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_48_3 dadda_fa_2_48_3/A dadda_fa_2_48_3/B dadda_fa_2_48_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/B dadda_fa_3_48_3/B sky130_fd_sc_hd__fa_1
XU$$3630 U$$4176/B1 U$$3674/A2 U$$4180/A1 U$$3674/B2 VGND VGND VPWR VPWR U$$3631/A
+ sky130_fd_sc_hd__a22o_1
XU$$4375 U$$4512/A1 U$$4381/A2 U$$4514/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4376/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4386 U$$4386/A VGND VGND VPWR VPWR U$$4386/Y sky130_fd_sc_hd__inv_1
XFILLER_77_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3641 U$$3641/A U$$3675/B VGND VGND VPWR VPWR U$$3641/X sky130_fd_sc_hd__xor2_1
XU$$3652 U$$3652/A1 U$$3664/A2 U$$3789/B1 U$$3664/B2 VGND VGND VPWR VPWR U$$3653/A
+ sky130_fd_sc_hd__a22o_1
XU$$4397 U$$4397/A U$$4397/B VGND VGND VPWR VPWR U$$4397/X sky130_fd_sc_hd__xor2_1
XFILLER_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3663 U$$3663/A U$$3663/B VGND VGND VPWR VPWR U$$3663/X sky130_fd_sc_hd__xor2_1
XFILLER_129_1209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3674 U$$3674/A1 U$$3674/A2 U$$4087/A1 U$$3674/B2 VGND VGND VPWR VPWR U$$3675/A
+ sky130_fd_sc_hd__a22o_1
XU$$2940 U$$2940/A U$$2972/B VGND VGND VPWR VPWR U$$2940/X sky130_fd_sc_hd__xor2_1
XFILLER_34_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_18_1 dadda_fa_5_18_1/A dadda_fa_5_18_1/B dadda_fa_5_18_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_19_0/B dadda_fa_7_18_0/A sky130_fd_sc_hd__fa_1
XU$$3685 U$$3685/A U$$3699/A VGND VGND VPWR VPWR U$$3685/X sky130_fd_sc_hd__xor2_1
XFILLER_52_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2951 U$$3088/A1 U$$2959/A2 U$$4186/A1 U$$2959/B2 VGND VGND VPWR VPWR U$$2952/A
+ sky130_fd_sc_hd__a22o_1
XU$$3696 U$$406/B1 U$$3696/A2 U$$3696/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3697/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2962 U$$2962/A U$$2966/B VGND VGND VPWR VPWR U$$2962/X sky130_fd_sc_hd__xor2_1
XU$$2973 U$$4480/A1 U$$2973/A2 U$$4482/A1 U$$2973/B2 VGND VGND VPWR VPWR U$$2974/A
+ sky130_fd_sc_hd__a22o_1
XU$$2984 U$$2984/A U$$3000/B VGND VGND VPWR VPWR U$$2984/X sky130_fd_sc_hd__xor2_1
XU$$2995 U$$3132/A1 U$$2997/A2 U$$3269/B1 U$$2997/B2 VGND VGND VPWR VPWR U$$2996/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_9_clk _442_/CLK VGND VGND VPWR VPWR _451_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_50_3 U$$1304/X U$$1437/X U$$1570/X VGND VGND VPWR VPWR dadda_fa_2_51_1/B
+ dadda_fa_2_50_4/B sky130_fd_sc_hd__fa_1
XU$$807 U$$944/A1 U$$809/A2 U$$944/B1 U$$809/B2 VGND VGND VPWR VPWR U$$808/A sky130_fd_sc_hd__a22o_1
XU$$818 U$$818/A U$$821/A VGND VGND VPWR VPWR U$$818/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_43_2 U$$891/X U$$1024/X U$$1157/X VGND VGND VPWR VPWR dadda_fa_2_44_3/B
+ dadda_fa_2_43_5/B sky130_fd_sc_hd__fa_1
XU$$829 U$$829/A U$$859/B VGND VGND VPWR VPWR U$$829/X sky130_fd_sc_hd__xor2_1
XFILLER_44_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_20_1 dadda_fa_4_20_1/A dadda_fa_4_20_1/B dadda_fa_4_20_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_21_0/B dadda_fa_5_20_1/B sky130_fd_sc_hd__fa_1
XFILLER_3_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_13_0 U$$33/X U$$166/X U$$299/X VGND VGND VPWR VPWR dadda_fa_5_14_0/A dadda_fa_5_13_1/A
+ sky130_fd_sc_hd__fa_1
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_803 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1707 U$$3157/B1 VGND VGND VPWR VPWR U$$2611/A1 sky130_fd_sc_hd__buf_6
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_65_3 dadda_fa_3_65_3/A dadda_fa_3_65_3/B dadda_fa_3_65_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_1/B dadda_fa_4_65_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_58_2 dadda_fa_3_58_2/A dadda_fa_3_58_2/B dadda_fa_3_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_1/A dadda_fa_4_58_2/B sky130_fd_sc_hd__fa_1
XFILLER_87_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_28_0 dadda_fa_6_28_0/A dadda_fa_6_28_0/B dadda_fa_6_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_29_0/B dadda_fa_7_28_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2203 U$$2203/A U$$2241/B VGND VGND VPWR VPWR U$$2203/X sky130_fd_sc_hd__xor2_1
XFILLER_35_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2214 U$$2625/A1 U$$2302/A2 U$$24/A1 U$$2302/B2 VGND VGND VPWR VPWR U$$2215/A sky130_fd_sc_hd__a22o_1
XFILLER_35_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2225 U$$2225/A U$$2269/B VGND VGND VPWR VPWR U$$2225/X sky130_fd_sc_hd__xor2_1
XU$$2236 U$$2508/B1 U$$2242/A2 U$$2375/A1 U$$2242/B2 VGND VGND VPWR VPWR U$$2237/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2247 U$$2247/A U$$2299/B VGND VGND VPWR VPWR U$$2247/X sky130_fd_sc_hd__xor2_1
XFILLER_90_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1502 U$$678/B1 U$$1374/X U$$545/A1 U$$1375/X VGND VGND VPWR VPWR U$$1503/A sky130_fd_sc_hd__a22o_1
XU$$2258 U$$3902/A1 U$$2274/A2 U$$66/B1 U$$2274/B2 VGND VGND VPWR VPWR U$$2259/A sky130_fd_sc_hd__a22o_1
XFILLER_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1513 U$$1513/A1 U$$1557/A2 U$$828/B1 U$$1557/B2 VGND VGND VPWR VPWR U$$1514/A
+ sky130_fd_sc_hd__a22o_1
XU$$1524 U$$1524/A U$$1554/B VGND VGND VPWR VPWR U$$1524/X sky130_fd_sc_hd__xor2_1
XFILLER_16_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2269 U$$2269/A U$$2269/B VGND VGND VPWR VPWR U$$2269/X sky130_fd_sc_hd__xor2_1
XU$$1535 U$$3042/A1 U$$1577/A2 U$$3042/B1 U$$1577/B2 VGND VGND VPWR VPWR U$$1536/A
+ sky130_fd_sc_hd__a22o_1
XU$$1546 U$$1546/A U$$1562/B VGND VGND VPWR VPWR U$$1546/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1557 U$$733/B1 U$$1557/A2 U$$600/A1 U$$1557/B2 VGND VGND VPWR VPWR U$$1558/A sky130_fd_sc_hd__a22o_1
XU$$1568 U$$1568/A U$$1588/B VGND VGND VPWR VPWR U$$1568/X sky130_fd_sc_hd__xor2_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_4__f_clk clkbuf_2_2_0_clk/X VGND VGND VPWR VPWR _634_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1579 U$$3221/B1 U$$1627/A2 U$$3088/A1 U$$1627/B2 VGND VGND VPWR VPWR U$$1580/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_777 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_229_ _353_/CLK _229_/D VGND VGND VPWR VPWR _229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_2 dadda_fa_2_60_2/A dadda_fa_2_60_2/B dadda_fa_2_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/A dadda_fa_3_60_3/A sky130_fd_sc_hd__fa_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater402 U$$809/A2 VGND VGND VPWR VPWR U$$765/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$209 final_adder.U$$703/A final_adder.U$$575/B1 final_adder.U$$209/B1
+ VGND VGND VPWR VPWR final_adder.U$$209/X sky130_fd_sc_hd__a21o_1
Xrepeater413 U$$668/A2 VGND VGND VPWR VPWR U$$622/A2 sky130_fd_sc_hd__buf_4
XFILLER_85_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater424 U$$457/A2 VGND VGND VPWR VPWR U$$447/A2 sky130_fd_sc_hd__buf_4
XFILLER_66_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_53_1 dadda_fa_2_53_1/A dadda_fa_2_53_1/B dadda_fa_2_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_0/CIN dadda_fa_3_53_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater435 U$$4114/X VGND VGND VPWR VPWR U$$4174/A2 sky130_fd_sc_hd__buf_6
Xrepeater446 U$$4/X VGND VGND VPWR VPWR U$$62/A2 sky130_fd_sc_hd__buf_2
XFILLER_38_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater457 U$$3910/A2 VGND VGND VPWR VPWR U$$3874/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_30_0 dadda_fa_5_30_0/A dadda_fa_5_30_0/B dadda_fa_5_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_31_0/A dadda_fa_6_30_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater468 U$$3805/A2 VGND VGND VPWR VPWR U$$3823/A2 sky130_fd_sc_hd__buf_8
XU$$4150 _568_/Q U$$4182/A2 _569_/Q U$$4182/B2 VGND VGND VPWR VPWR U$$4151/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_46_0 U$$2759/X U$$2892/X U$$3025/X VGND VGND VPWR VPWR dadda_fa_3_47_0/B
+ dadda_fa_3_46_2/B sky130_fd_sc_hd__fa_1
XFILLER_93_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater479 U$$3429/X VGND VGND VPWR VPWR U$$3497/A2 sky130_fd_sc_hd__buf_6
XU$$4161 U$$4161/A U$$4175/B VGND VGND VPWR VPWR U$$4161/X sky130_fd_sc_hd__xor2_1
XFILLER_26_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4172 U$$4444/B1 U$$4174/A2 U$$4446/B1 U$$4174/B2 VGND VGND VPWR VPWR U$$4173/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4183 U$$4183/A U$$4183/B VGND VGND VPWR VPWR U$$4183/X sky130_fd_sc_hd__xor2_1
XFILLER_81_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4194 U$$4468/A1 U$$4196/A2 U$$4194/B1 U$$4196/B2 VGND VGND VPWR VPWR U$$4195/A
+ sky130_fd_sc_hd__a22o_1
XU$$3460 U$$3460/A U$$3561/A VGND VGND VPWR VPWR U$$3460/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3471 U$$4293/A1 U$$3545/A2 U$$4158/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3472/A
+ sky130_fd_sc_hd__a22o_1
XU$$3482 U$$3482/A U$$3490/B VGND VGND VPWR VPWR U$$3482/X sky130_fd_sc_hd__xor2_1
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3493 U$$3493/A1 U$$3497/A2 U$$3495/A1 U$$3497/B2 VGND VGND VPWR VPWR U$$3494/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2770 U$$3042/B1 U$$2814/A2 U$$2909/A1 U$$2814/B2 VGND VGND VPWR VPWR U$$2771/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2781 U$$2781/A U$$2813/B VGND VGND VPWR VPWR U$$2781/X sky130_fd_sc_hd__xor2_1
XFILLER_209_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2792 U$$463/A1 U$$2798/A2 U$$463/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2793/A sky130_fd_sc_hd__a22o_1
XFILLER_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_75_2 dadda_fa_4_75_2/A dadda_fa_4_75_2/B dadda_fa_4_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/CIN dadda_fa_5_75_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_68_1 dadda_fa_4_68_1/A dadda_fa_4_68_1/B dadda_fa_4_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/B dadda_fa_5_68_1/B sky130_fd_sc_hd__fa_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput205 c[53] VGND VGND VPWR VPWR input205/X sky130_fd_sc_hd__clkbuf_4
Xinput216 c[63] VGND VGND VPWR VPWR input216/X sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_7_45_0 dadda_fa_7_45_0/A dadda_fa_7_45_0/B dadda_fa_7_45_0/CIN VGND VGND
+ VPWR VPWR _470_/D _341_/D sky130_fd_sc_hd__fa_1
Xinput227 c[73] VGND VGND VPWR VPWR input227/X sky130_fd_sc_hd__clkbuf_4
XTAP_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput238 c[83] VGND VGND VPWR VPWR input238/X sky130_fd_sc_hd__buf_2
XFILLER_102_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_1_35_0 U$$77/X U$$210/X VGND VGND VPWR VPWR dadda_fa_2_36_5/B dadda_fa_3_35_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_130_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$710 final_adder.U$$710/A final_adder.U$$710/B VGND VGND VPWR VPWR
+ _256_/D sky130_fd_sc_hd__xor2_1
Xinput249 c[93] VGND VGND VPWR VPWR input249/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$721 final_adder.U$$721/A final_adder.U$$721/B VGND VGND VPWR VPWR
+ _267_/D sky130_fd_sc_hd__xor2_1
XTAP_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_691 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$732 final_adder.U$$732/A final_adder.U$$732/B VGND VGND VPWR VPWR
+ _278_/D sky130_fd_sc_hd__xor2_4
XTAP_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$743 final_adder.U$$743/A final_adder.U$$743/B VGND VGND VPWR VPWR
+ _289_/D sky130_fd_sc_hd__xor2_4
XFILLER_57_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$604 U$$878/A1 U$$616/A2 U$$880/A1 U$$616/B2 VGND VGND VPWR VPWR U$$605/A sky130_fd_sc_hd__a22o_1
XFILLER_1_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_580_ _582_/CLK _580_/D VGND VGND VPWR VPWR _580_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater980 U$$3286/B VGND VGND VPWR VPWR U$$3236/B sky130_fd_sc_hd__buf_8
XFILLER_84_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$615 U$$615/A U$$659/B VGND VGND VPWR VPWR U$$615/X sky130_fd_sc_hd__xor2_1
XU$$626 U$$761/B1 U$$632/A2 U$$628/A1 U$$632/B2 VGND VGND VPWR VPWR U$$627/A sky130_fd_sc_hd__a22o_1
XFILLER_57_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater991 U$$3145/B VGND VGND VPWR VPWR U$$3121/B sky130_fd_sc_hd__buf_6
XU$$637 U$$637/A U$$651/B VGND VGND VPWR VPWR U$$637/X sky130_fd_sc_hd__xor2_1
XFILLER_16_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$648 U$$648/A1 U$$650/A2 U$$648/B1 U$$650/B2 VGND VGND VPWR VPWR U$$649/A sky130_fd_sc_hd__a22o_1
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$659 U$$659/A U$$659/B VGND VGND VPWR VPWR U$$659/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_731 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1504 U$$3346/A1 VGND VGND VPWR VPWR U$$467/B1 sky130_fd_sc_hd__buf_6
Xrepeater1515 _576_/Q VGND VGND VPWR VPWR U$$4440/A1 sky130_fd_sc_hd__buf_8
XFILLER_125_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1526 U$$52/A1 VGND VGND VPWR VPWR U$$874/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1537 U$$3475/A1 VGND VGND VPWR VPWR U$$50/A1 sky130_fd_sc_hd__buf_8
Xrepeater1548 U$$4154/B1 VGND VGND VPWR VPWR U$$2375/A1 sky130_fd_sc_hd__buf_4
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1559 U$$3741/B1 VGND VGND VPWR VPWR U$$3056/B1 sky130_fd_sc_hd__buf_4
XFILLER_180_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_70_1 dadda_fa_3_70_1/A dadda_fa_3_70_1/B dadda_fa_3_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_0/CIN dadda_fa_4_70_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_63_0 dadda_fa_3_63_0/A dadda_fa_3_63_0/B dadda_fa_3_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_0/B dadda_fa_4_63_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2000 U$$3505/B1 U$$1922/X U$$3372/A1 U$$1923/X VGND VGND VPWR VPWR U$$2001/A sky130_fd_sc_hd__a22o_1
XFILLER_208_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2011 U$$2011/A U$$2011/B VGND VGND VPWR VPWR U$$2011/X sky130_fd_sc_hd__xor2_1
XU$$2022 U$$3253/B1 U$$2028/A2 U$$3255/B1 U$$2028/B2 VGND VGND VPWR VPWR U$$2023/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2033 U$$2033/A U$$2039/B VGND VGND VPWR VPWR U$$2033/X sky130_fd_sc_hd__xor2_1
XFILLER_90_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2044 U$$946/B1 U$$2052/A2 U$$2318/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2045/A
+ sky130_fd_sc_hd__a22o_1
XU$$1310 U$$1310/A U$$1310/B VGND VGND VPWR VPWR U$$1310/X sky130_fd_sc_hd__xor2_1
XFILLER_16_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2055 _645_/Q VGND VGND VPWR VPWR U$$2055/Y sky130_fd_sc_hd__inv_1
XU$$1321 U$$634/B1 U$$1355/A2 U$$501/A1 U$$1355/B2 VGND VGND VPWR VPWR U$$1322/A sky130_fd_sc_hd__a22o_1
XU$$2066 U$$2066/A U$$2110/B VGND VGND VPWR VPWR U$$2066/X sky130_fd_sc_hd__xor2_1
XU$$2077 U$$20/B1 U$$2115/A2 U$$2077/B1 U$$2115/B2 VGND VGND VPWR VPWR U$$2078/A sky130_fd_sc_hd__a22o_1
XU$$1332 U$$1332/A U$$1332/B VGND VGND VPWR VPWR U$$1332/X sky130_fd_sc_hd__xor2_1
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2088 U$$2088/A U$$2130/B VGND VGND VPWR VPWR U$$2088/X sky130_fd_sc_hd__xor2_1
XU$$1343 U$$2848/B1 U$$1345/A2 U$$658/B1 U$$1345/B2 VGND VGND VPWR VPWR U$$1344/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1354 U$$1354/A U$$1356/B VGND VGND VPWR VPWR U$$1354/X sky130_fd_sc_hd__xor2_1
XFILLER_210_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2099 U$$44/A1 U$$2115/A2 U$$46/A1 U$$2115/B2 VGND VGND VPWR VPWR U$$2100/A sky130_fd_sc_hd__a22o_1
XU$$1365 U$$817/A1 U$$1367/A2 U$$817/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1366/A sky130_fd_sc_hd__a22o_1
XU$$1376 U$$1376/A1 U$$1428/A2 U$$8/A1 U$$1428/B2 VGND VGND VPWR VPWR U$$1377/A sky130_fd_sc_hd__a22o_1
XU$$1387 U$$1387/A U$$1425/B VGND VGND VPWR VPWR U$$1387/X sky130_fd_sc_hd__xor2_1
XFILLER_176_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_120_0 dadda_fa_7_120_0/A dadda_fa_7_120_0/B dadda_fa_7_120_0/CIN VGND
+ VGND VPWR VPWR _545_/D _416_/D sky130_fd_sc_hd__fa_1
XU$$1398 U$$987/A1 U$$1424/A2 U$$2494/B1 U$$1424/B2 VGND VGND VPWR VPWR U$$1399/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_85_1 dadda_fa_5_85_1/A dadda_fa_5_85_1/B dadda_fa_5_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_86_0/B dadda_fa_7_85_0/A sky130_fd_sc_hd__fa_2
XFILLER_7_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_78_0 dadda_fa_5_78_0/A dadda_fa_5_78_0/B dadda_fa_5_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_79_0/A dadda_fa_6_78_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_144_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_77_8 input231/X dadda_fa_1_77_8/B dadda_fa_1_77_8/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_78_3/A dadda_fa_3_77_0/A sky130_fd_sc_hd__fa_2
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1087 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$50 _474_/Q _346_/Q VGND VGND VPWR VPWR final_adder.U$$545/B1 final_adder.U$$672/A
+ sky130_fd_sc_hd__ha_1
XFILLER_199_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$61 _485_/Q _357_/Q VGND VGND VPWR VPWR final_adder.U$$189/B1 final_adder.U$$683/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3290 U$$3423/B VGND VGND VPWR VPWR U$$3290/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$72 _496_/Q _368_/Q VGND VGND VPWR VPWR final_adder.U$$567/B1 final_adder.U$$694/A
+ sky130_fd_sc_hd__ha_1
XFILLER_53_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$83 _507_/Q _379_/Q VGND VGND VPWR VPWR final_adder.U$$211/B1 final_adder.U$$705/A
+ sky130_fd_sc_hd__ha_1
XFILLER_198_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$94 _518_/Q _390_/Q VGND VGND VPWR VPWR final_adder.U$$589/B1 final_adder.U$$716/A
+ sky130_fd_sc_hd__ha_1
XFILLER_55_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_471 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_80_0 dadda_fa_4_80_0/A dadda_fa_4_80_0/B dadda_fa_4_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/A dadda_fa_5_80_1/A sky130_fd_sc_hd__fa_1
XFILLER_162_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_101_3 dadda_fa_3_101_3/A dadda_fa_3_101_3/B dadda_fa_3_101_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_102_1/B dadda_fa_4_101_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$551 final_adder.U$$678/A final_adder.U$$678/B final_adder.U$$551/B1
+ VGND VGND VPWR VPWR final_adder.U$$679/B sky130_fd_sc_hd__a21o_1
XTAP_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_632_ _633_/CLK _632_/D VGND VGND VPWR VPWR _632_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$401 U$$401/A U$$411/A VGND VGND VPWR VPWR U$$401/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_108_0 dadda_fa_6_108_0/A dadda_fa_6_108_0/B dadda_fa_6_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_109_0/B dadda_fa_7_108_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$573 final_adder.U$$700/A final_adder.U$$700/B final_adder.U$$573/B1
+ VGND VGND VPWR VPWR final_adder.U$$701/B sky130_fd_sc_hd__a21o_1
XTAP_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$412 _622_/Q VGND VGND VPWR VPWR U$$414/B sky130_fd_sc_hd__inv_1
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$423 U$$695/B1 U$$447/A2 U$$562/A1 U$$447/B2 VGND VGND VPWR VPWR U$$424/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$595 final_adder.U$$722/A final_adder.U$$722/B final_adder.U$$595/B1
+ VGND VGND VPWR VPWR final_adder.U$$723/B sky130_fd_sc_hd__a21o_1
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$434 U$$434/A U$$456/B VGND VGND VPWR VPWR U$$434/X sky130_fd_sc_hd__xor2_1
XFILLER_44_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_563_ _569_/CLK _563_/D VGND VGND VPWR VPWR _563_/Q sky130_fd_sc_hd__dfxtp_4
XU$$445 U$$582/A1 U$$447/A2 U$$582/B1 U$$447/B2 VGND VGND VPWR VPWR U$$446/A sky130_fd_sc_hd__a22o_1
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$456 U$$456/A U$$456/B VGND VGND VPWR VPWR U$$456/X sky130_fd_sc_hd__xor2_1
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_28_3 dadda_fa_3_28_3/A dadda_fa_3_28_3/B dadda_fa_3_28_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_29_1/B dadda_fa_4_28_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_72_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$467 U$$467/A1 U$$499/A2 U$$467/B1 U$$499/B2 VGND VGND VPWR VPWR U$$468/A sky130_fd_sc_hd__a22o_1
XU$$478 U$$478/A U$$484/B VGND VGND VPWR VPWR U$$478/X sky130_fd_sc_hd__xor2_1
XU$$489 U$$624/B1 U$$491/A2 U$$491/A1 U$$491/B2 VGND VGND VPWR VPWR U$$490/A sky130_fd_sc_hd__a22o_1
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_494_ _494_/CLK _494_/D VGND VGND VPWR VPWR _494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_95_0 dadda_fa_6_95_0/A dadda_fa_6_95_0/B dadda_fa_6_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_96_0/B dadda_fa_7_95_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_139_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1301 U$$4490/B1 VGND VGND VPWR VPWR U$$930/A1 sky130_fd_sc_hd__buf_4
Xrepeater1312 U$$3805/A1 VGND VGND VPWR VPWR U$$3942/A1 sky130_fd_sc_hd__buf_4
XFILLER_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1323 U$$3799/B1 VGND VGND VPWR VPWR U$$924/A1 sky130_fd_sc_hd__buf_6
XFILLER_158_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1334 U$$3934/B1 VGND VGND VPWR VPWR U$$922/A1 sky130_fd_sc_hd__buf_6
XFILLER_158_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1345 U$$4206/B1 VGND VGND VPWR VPWR U$$918/B1 sky130_fd_sc_hd__buf_6
XFILLER_119_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1356 U$$3791/B1 VGND VGND VPWR VPWR U$$916/A1 sky130_fd_sc_hd__buf_4
XFILLER_180_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1367 _594_/Q VGND VGND VPWR VPWR U$$3789/B1 sky130_fd_sc_hd__buf_4
Xrepeater1378 _593_/Q VGND VGND VPWR VPWR U$$4198/B1 sky130_fd_sc_hd__buf_6
Xrepeater1389 U$$3783/B1 VGND VGND VPWR VPWR U$$2415/A1 sky130_fd_sc_hd__buf_6
XFILLER_79_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_30_3 U$$1264/X U$$1397/X U$$1530/X VGND VGND VPWR VPWR dadda_fa_3_31_2/A
+ dadda_fa_3_30_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_91_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$990 U$$990/A U$$994/B VGND VGND VPWR VPWR U$$990/X sky130_fd_sc_hd__xor2_1
XFILLER_51_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1140 U$$2508/B1 U$$1146/A2 U$$2375/A1 U$$1146/B2 VGND VGND VPWR VPWR U$$1141/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1151 U$$1151/A U$$1151/B VGND VGND VPWR VPWR U$$1151/X sky130_fd_sc_hd__xor2_1
XU$$1162 U$$749/B1 U$$1190/A2 U$$68/A1 U$$1190/B2 VGND VGND VPWR VPWR U$$1163/A sky130_fd_sc_hd__a22o_1
XU$$1173 U$$1173/A U$$1177/B VGND VGND VPWR VPWR U$$1173/X sky130_fd_sc_hd__xor2_1
XFILLER_210_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1184 U$$634/B1 U$$1224/A2 U$$501/A1 U$$1224/B2 VGND VGND VPWR VPWR U$$1185/A sky130_fd_sc_hd__a22o_1
XU$$1195 U$$1195/A U$$1195/B VGND VGND VPWR VPWR U$$1195/X sky130_fd_sc_hd__xor2_1
XFILLER_31_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_82_6 U$$3629/X U$$3762/X U$$3895/X VGND VGND VPWR VPWR dadda_fa_2_83_3/B
+ dadda_fa_2_82_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_75_5 U$$3615/X U$$3748/X U$$3881/X VGND VGND VPWR VPWR dadda_fa_2_76_2/A
+ dadda_fa_2_75_5/A sky130_fd_sc_hd__fa_1
XFILLER_86_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_4 U$$4133/X U$$4266/X U$$4399/X VGND VGND VPWR VPWR dadda_fa_2_69_1/CIN
+ dadda_fa_2_68_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1010 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_2 dadda_fa_4_38_2/A dadda_fa_4_38_2/B dadda_fa_4_38_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/CIN dadda_fa_5_38_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _179_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_129 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_599 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_3 U$$1330/X U$$1463/X U$$1596/X VGND VGND VPWR VPWR dadda_fa_1_64_6/B
+ dadda_fa_1_63_8/B sky130_fd_sc_hd__fa_1
XTAP_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_40_2 dadda_fa_3_40_2/A dadda_fa_3_40_2/B dadda_fa_3_40_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_1/A dadda_fa_4_40_2/B sky130_fd_sc_hd__fa_1
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$370 final_adder.U$$370/A final_adder.U$$370/B VGND VGND VPWR VPWR
+ final_adder.U$$370/X sky130_fd_sc_hd__and2_1
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_615_ _615_/CLK _615_/D VGND VGND VPWR VPWR _615_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_205_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_33_1 dadda_fa_3_33_1/A dadda_fa_3_33_1/B dadda_fa_3_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_0/CIN dadda_fa_4_33_2/A sky130_fd_sc_hd__fa_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$220 U$$220/A U$$226/B VGND VGND VPWR VPWR U$$220/X sky130_fd_sc_hd__xor2_1
XFILLER_205_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$231 U$$368/A1 U$$259/A2 U$$96/A1 U$$259/B2 VGND VGND VPWR VPWR U$$232/A sky130_fd_sc_hd__a22o_1
XU$$242 U$$242/A U$$250/B VGND VGND VPWR VPWR U$$242/X sky130_fd_sc_hd__xor2_1
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_10_0 dadda_fa_6_10_0/A dadda_fa_6_10_0/B dadda_fa_6_10_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_11_0/B dadda_fa_7_10_0/CIN sky130_fd_sc_hd__fa_1
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_26_0 U$$1123/X U$$1256/X U$$1389/X VGND VGND VPWR VPWR dadda_fa_4_27_0/B
+ dadda_fa_4_26_1/CIN sky130_fd_sc_hd__fa_1
XU$$253 U$$527/A1 U$$259/A2 U$$253/B1 U$$259/B2 VGND VGND VPWR VPWR U$$254/A sky130_fd_sc_hd__a22o_1
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$264 U$$264/A U$$264/B VGND VGND VPWR VPWR U$$264/X sky130_fd_sc_hd__xor2_1
XFILLER_60_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_546_ _547_/CLK _546_/D VGND VGND VPWR VPWR _546_/Q sky130_fd_sc_hd__dfxtp_1
XU$$275 _620_/Q VGND VGND VPWR VPWR U$$277/B sky130_fd_sc_hd__inv_1
XFILLER_75_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$286 U$$12/A1 U$$318/A2 U$$14/A1 U$$318/B2 VGND VGND VPWR VPWR U$$287/A sky130_fd_sc_hd__a22o_1
XFILLER_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$297 U$$297/A U$$309/B VGND VGND VPWR VPWR U$$297/X sky130_fd_sc_hd__xor2_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_477_ _478_/CLK _477_/D VGND VGND VPWR VPWR _477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3 U$$3/A U$$3/B VGND VGND VPWR VPWR U$$3/X sky130_fd_sc_hd__and2_1
XFILLER_12_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput306 _197_/Q VGND VGND VPWR VPWR o[29] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_5 dadda_fa_2_92_5/A dadda_fa_2_92_5/B dadda_fa_2_92_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_93_2/A dadda_fa_4_92_0/A sky130_fd_sc_hd__fa_1
Xrepeater1120 U$$996/B VGND VGND VPWR VPWR U$$994/B sky130_fd_sc_hd__buf_6
Xoutput317 _207_/Q VGND VGND VPWR VPWR o[39] sky130_fd_sc_hd__buf_2
Xrepeater1131 U$$897/B VGND VGND VPWR VPWR U$$879/B sky130_fd_sc_hd__buf_6
Xoutput328 _217_/Q VGND VGND VPWR VPWR o[49] sky130_fd_sc_hd__buf_2
XFILLER_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1142 U$$810/B VGND VGND VPWR VPWR U$$766/B sky130_fd_sc_hd__buf_6
Xrepeater1153 U$$669/B VGND VGND VPWR VPWR U$$665/B sky130_fd_sc_hd__buf_6
Xoutput339 _227_/Q VGND VGND VPWR VPWR o[59] sky130_fd_sc_hd__buf_2
XFILLER_141_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_85_4 dadda_fa_2_85_4/A dadda_fa_2_85_4/B dadda_fa_2_85_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/CIN dadda_fa_3_85_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1164 U$$309/B VGND VGND VPWR VPWR U$$319/B sky130_fd_sc_hd__buf_6
XFILLER_113_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1175 U$$264/B VGND VGND VPWR VPWR U$$226/B sky130_fd_sc_hd__buf_6
XFILLER_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1186 U$$85/B VGND VGND VPWR VPWR U$$81/B sky130_fd_sc_hd__buf_6
XFILLER_142_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1197 U$$2872/B1 VGND VGND VPWR VPWR U$$3285/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_78_3 dadda_fa_2_78_3/A dadda_fa_2_78_3/B dadda_fa_2_78_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/B dadda_fa_3_78_3/B sky130_fd_sc_hd__fa_1
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_48_1 dadda_fa_5_48_1/A dadda_fa_5_48_1/B dadda_fa_5_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_49_0/B dadda_fa_7_48_0/A sky130_fd_sc_hd__fa_1
XFILLER_82_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_101_2 U$$3401/X U$$3534/X U$$3667/X VGND VGND VPWR VPWR dadda_fa_3_102_2/B
+ dadda_fa_3_101_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_122_1 input154/X dadda_fa_5_122_1/B dadda_ha_4_122_0/SUM VGND VGND VPWR
+ VPWR dadda_fa_6_123_0/B dadda_fa_7_122_0/A sky130_fd_sc_hd__fa_1
XFILLER_177_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_115_0 dadda_fa_5_115_0/A dadda_fa_5_115_0/B dadda_fa_5_115_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_116_0/A dadda_fa_6_115_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_80_3 U$$2295/X U$$2428/X U$$2561/X VGND VGND VPWR VPWR dadda_fa_2_81_1/CIN
+ dadda_fa_2_80_4/B sky130_fd_sc_hd__fa_1
XFILLER_104_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_73_2 U$$2680/X U$$2813/X U$$2946/X VGND VGND VPWR VPWR dadda_fa_2_74_1/A
+ dadda_fa_2_73_4/A sky130_fd_sc_hd__fa_1
XFILLER_24_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_50_1 dadda_fa_4_50_1/A dadda_fa_4_50_1/B dadda_fa_4_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/B dadda_fa_5_50_1/B sky130_fd_sc_hd__fa_1
XFILLER_115_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_66_1 U$$2932/X U$$3065/X U$$3198/X VGND VGND VPWR VPWR dadda_fa_2_67_0/CIN
+ dadda_fa_2_66_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_2_100_4 U$$4064/X U$$4197/X VGND VGND VPWR VPWR dadda_fa_3_101_2/CIN dadda_fa_4_100_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_101_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_43_0 dadda_fa_4_43_0/A dadda_fa_4_43_0/B dadda_fa_4_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/A dadda_fa_5_43_1/A sky130_fd_sc_hd__fa_1
XFILLER_98_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_59_0 U$$1588/X U$$1721/X U$$1854/X VGND VGND VPWR VPWR dadda_fa_2_60_0/B
+ dadda_fa_2_59_3/B sky130_fd_sc_hd__fa_1
XFILLER_111_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_439 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_400_ _566_/CLK _400_/D VGND VGND VPWR VPWR _400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1909 U$$2318/B1 U$$1909/A2 U$$3418/A1 U$$1909/B2 VGND VGND VPWR VPWR U$$1910/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_612 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_331_ _463_/CLK _331_/D VGND VGND VPWR VPWR _331_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_262_ _520_/CLK _262_/D VGND VGND VPWR VPWR _262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_193_ _207_/CLK _193_/D VGND VGND VPWR VPWR _193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_95_3 dadda_fa_3_95_3/A dadda_fa_3_95_3/B dadda_fa_3_95_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_1/B dadda_fa_4_95_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_506 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_88_2 dadda_fa_3_88_2/A dadda_fa_3_88_2/B dadda_fa_3_88_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_1/A dadda_fa_4_88_2/B sky130_fd_sc_hd__fa_1
XFILLER_150_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_55_1 U$$516/X U$$649/X VGND VGND VPWR VPWR dadda_fa_1_56_8/A dadda_fa_2_55_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_58_0 dadda_fa_6_58_0/A dadda_fa_6_58_0/B dadda_fa_6_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_59_0/B dadda_fa_7_58_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater809 U$$2302/B2 VGND VGND VPWR VPWR U$$2248/B2 sky130_fd_sc_hd__buf_6
XU$$4502 U$$4502/A1 U$$4388/X U$$4504/A1 U$$4389/X VGND VGND VPWR VPWR U$$4503/A sky130_fd_sc_hd__a22o_1
XFILLER_110_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4513 U$$4513/A U$$4513/B VGND VGND VPWR VPWR U$$4513/X sky130_fd_sc_hd__xor2_1
XFILLER_2_46 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_61_0 U$$129/X U$$262/X U$$395/X VGND VGND VPWR VPWR dadda_fa_1_62_5/CIN
+ dadda_fa_1_61_7/CIN sky130_fd_sc_hd__fa_1
XU$$16 U$$16/A1 U$$8/A2 U$$18/A1 U$$8/B2 VGND VGND VPWR VPWR U$$17/A sky130_fd_sc_hd__a22o_1
XU$$3801 U$$4075/A1 U$$3805/A2 U$$3803/A1 U$$3805/B2 VGND VGND VPWR VPWR U$$3802/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3812 U$$3812/A U$$3816/B VGND VGND VPWR VPWR U$$3812/X sky130_fd_sc_hd__xor2_1
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_117_2 U$$4497/X input148/X dadda_fa_4_117_2/CIN VGND VGND VPWR VPWR dadda_fa_5_118_0/CIN
+ dadda_fa_5_117_1/CIN sky130_fd_sc_hd__fa_1
XU$$3823 U$$4369/B1 U$$3823/A2 U$$4236/A1 U$$3823/B2 VGND VGND VPWR VPWR U$$3824/A
+ sky130_fd_sc_hd__a22o_1
XU$$27 U$$27/A U$$57/B VGND VGND VPWR VPWR U$$27/X sky130_fd_sc_hd__xor2_1
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$38 U$$38/A1 U$$62/A2 U$$40/A1 U$$62/B2 VGND VGND VPWR VPWR U$$39/A sky130_fd_sc_hd__a22o_1
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$49 U$$49/A U$$85/B VGND VGND VPWR VPWR U$$49/X sky130_fd_sc_hd__xor2_1
XU$$3834 U$$3834/A U$$3835/A VGND VGND VPWR VPWR U$$3834/X sky130_fd_sc_hd__xor2_1
XU$$3845 U$$3845/A U$$3895/B VGND VGND VPWR VPWR U$$3845/X sky130_fd_sc_hd__xor2_1
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3856 U$$4402/B1 U$$3970/A2 U$$4269/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3857/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3867 U$$3867/A U$$3949/B VGND VGND VPWR VPWR U$$3867/X sky130_fd_sc_hd__xor2_1
XU$$3878 _569_/Q U$$3916/A2 U$$4154/A1 U$$3916/B2 VGND VGND VPWR VPWR U$$3879/A sky130_fd_sc_hd__a22o_1
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3889 U$$3889/A U$$3917/B VGND VGND VPWR VPWR U$$3889/X sky130_fd_sc_hd__xor2_1
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_529_ _566_/CLK _529_/D VGND VGND VPWR VPWR _529_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_18 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_330 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_29 _282_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4395_1776 VGND VGND VPWR VPWR U$$4395_1776/HI U$$4395/B sky130_fd_sc_hd__conb_1
XFILLER_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_90_2 U$$4044/X U$$4177/X U$$4310/X VGND VGND VPWR VPWR dadda_fa_3_91_1/A
+ dadda_fa_3_90_3/A sky130_fd_sc_hd__fa_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_83_1 input238/X dadda_fa_2_83_1/B dadda_fa_2_83_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_84_0/CIN dadda_fa_3_83_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_60_0 dadda_fa_5_60_0/A dadda_fa_5_60_0/B dadda_fa_5_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_61_0/A dadda_fa_6_60_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_76_0 dadda_fa_2_76_0/A dadda_fa_2_76_0/B dadda_fa_2_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_0/B dadda_fa_3_76_2/B sky130_fd_sc_hd__fa_1
XFILLER_130_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_52_7 U$$3170/X U$$3303/X U$$3436/X VGND VGND VPWR VPWR dadda_fa_2_53_2/CIN
+ dadda_fa_2_52_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_98_1 dadda_fa_4_98_1/A dadda_fa_4_98_1/B dadda_fa_4_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/B dadda_fa_5_98_1/B sky130_fd_sc_hd__fa_1
XFILLER_30_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_75_0 dadda_fa_7_75_0/A dadda_fa_7_75_0/B dadda_fa_7_75_0/CIN VGND VGND
+ VPWR VPWR _500_/D _371_/D sky130_fd_sc_hd__fa_1
XFILLER_127_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_274 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3108 U$$4478/A1 U$$3144/A2 U$$4480/A1 U$$3144/B2 VGND VGND VPWR VPWR U$$3109/A
+ sky130_fd_sc_hd__a22o_1
XU$$3119 U$$3119/A U$$3121/B VGND VGND VPWR VPWR U$$3119/X sky130_fd_sc_hd__xor2_1
XFILLER_86_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2407 U$$3503/A1 U$$2437/A2 U$$628/A1 U$$2437/B2 VGND VGND VPWR VPWR U$$2408/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2418 U$$2418/A U$$2418/B VGND VGND VPWR VPWR U$$2418/X sky130_fd_sc_hd__xor2_1
XFILLER_36_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2429 U$$3934/B1 U$$2451/A2 U$$785/B1 U$$2451/B2 VGND VGND VPWR VPWR U$$2430/A
+ sky130_fd_sc_hd__a22o_1
XU$$1706 U$$1843/A1 U$$1710/A2 U$$3352/A1 U$$1710/B2 VGND VGND VPWR VPWR U$$1707/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1717 U$$1717/A U$$1719/B VGND VGND VPWR VPWR U$$1717/X sky130_fd_sc_hd__xor2_1
XFILLER_36_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1728 U$$358/A1 U$$1736/A2 U$$86/A1 U$$1736/B2 VGND VGND VPWR VPWR U$$1729/A sky130_fd_sc_hd__a22o_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1739 U$$1739/A U$$1747/B VGND VGND VPWR VPWR U$$1739/X sky130_fd_sc_hd__xor2_1
XFILLER_54_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_314_ _441_/CLK _314_/D VGND VGND VPWR VPWR _314_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_245_ _372_/CLK _245_/D VGND VGND VPWR VPWR _245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1083 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput16 a[23] VGND VGND VPWR VPWR _639_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput27 a[33] VGND VGND VPWR VPWR _649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput38 a[43] VGND VGND VPWR VPWR _659_/D sky130_fd_sc_hd__clkbuf_1
X_176_ _428_/CLK _176_/D VGND VGND VPWR VPWR _176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput49 a[53] VGND VGND VPWR VPWR _669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_182_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_93_0 dadda_fa_3_93_0/A dadda_fa_3_93_0/B dadda_fa_3_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_0/B dadda_fa_4_93_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_202_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater606 U$$1511/X VGND VGND VPWR VPWR U$$1635/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_172_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater617 U$$1474/A2 VGND VGND VPWR VPWR U$$1458/A2 sky130_fd_sc_hd__buf_4
XFILLER_81_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater628 U$$1237/X VGND VGND VPWR VPWR U$$1323/A2 sky130_fd_sc_hd__buf_4
XFILLER_77_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4310 U$$4310/A _679_/Q VGND VGND VPWR VPWR U$$4310/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_55_5 dadda_fa_2_55_5/A dadda_fa_2_55_5/B dadda_fa_2_55_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_2/A dadda_fa_4_55_0/A sky130_fd_sc_hd__fa_2
XU$$4321 _585_/Q U$$4335/A2 _586_/Q U$$4333/B2 VGND VGND VPWR VPWR U$$4322/A sky130_fd_sc_hd__a22o_1
Xrepeater639 U$$1100/X VGND VGND VPWR VPWR U$$1208/A2 sky130_fd_sc_hd__buf_6
XFILLER_120_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4332 U$$4332/A U$$4334/B VGND VGND VPWR VPWR U$$4332/X sky130_fd_sc_hd__xor2_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4343 U$$4480/A1 U$$4251/X U$$4482/A1 U$$4345/B2 VGND VGND VPWR VPWR U$$4344/A
+ sky130_fd_sc_hd__a22o_1
XU$$4354 U$$4354/A U$$4382/B VGND VGND VPWR VPWR U$$4354/X sky130_fd_sc_hd__xor2_1
XU$$3620 _577_/Q U$$3664/A2 _578_/Q U$$3664/B2 VGND VGND VPWR VPWR U$$3621/A sky130_fd_sc_hd__a22o_1
XU$$4365 U$$4500/B1 U$$4369/A2 U$$805/A1 U$$4369/B2 VGND VGND VPWR VPWR U$$4366/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_48_4 dadda_fa_2_48_4/A dadda_fa_2_48_4/B dadda_fa_2_48_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/CIN dadda_fa_3_48_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4376 U$$4376/A U$$4383/A VGND VGND VPWR VPWR U$$4376/X sky130_fd_sc_hd__xor2_1
XU$$3631 U$$3631/A U$$3675/B VGND VGND VPWR VPWR U$$3631/X sky130_fd_sc_hd__xor2_1
XFILLER_203_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4387 U$$4387/A U$$4387/B VGND VGND VPWR VPWR U$$4387/X sky130_fd_sc_hd__and2_1
XU$$3642 U$$3642/A1 U$$3674/A2 U$$3779/B1 U$$3674/B2 VGND VGND VPWR VPWR U$$3643/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3653 U$$3653/A U$$3663/B VGND VGND VPWR VPWR U$$3653/X sky130_fd_sc_hd__xor2_1
XU$$4398 _555_/Q U$$4388/X _556_/Q U$$4438/B2 VGND VGND VPWR VPWR U$$4399/A sky130_fd_sc_hd__a22o_1
XFILLER_53_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3664 U$$4075/A1 U$$3664/A2 U$$3803/A1 U$$3664/B2 VGND VGND VPWR VPWR U$$3665/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2930 U$$2930/A U$$2972/B VGND VGND VPWR VPWR U$$2930/X sky130_fd_sc_hd__xor2_1
XU$$3675 U$$3675/A U$$3675/B VGND VGND VPWR VPWR U$$3675/X sky130_fd_sc_hd__xor2_1
XU$$3686 U$$4508/A1 U$$3688/A2 U$$4510/A1 U$$3688/B2 VGND VGND VPWR VPWR U$$3687/A
+ sky130_fd_sc_hd__a22o_1
XU$$2941 U$$201/A1 U$$2943/A2 U$$3626/B1 U$$2943/B2 VGND VGND VPWR VPWR U$$2942/A
+ sky130_fd_sc_hd__a22o_1
XU$$2952 U$$2952/A U$$2988/B VGND VGND VPWR VPWR U$$2952/X sky130_fd_sc_hd__xor2_1
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3697 U$$3697/A U$$3698/A VGND VGND VPWR VPWR U$$3697/X sky130_fd_sc_hd__xor2_1
XFILLER_93_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2963 U$$3783/B1 U$$2981/A2 U$$2963/B1 U$$2981/B2 VGND VGND VPWR VPWR U$$2964/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2974 U$$2974/A U$$3008/B VGND VGND VPWR VPWR U$$2974/X sky130_fd_sc_hd__xor2_1
XU$$2985 U$$3122/A1 U$$2997/A2 U$$3124/A1 U$$2997/B2 VGND VGND VPWR VPWR U$$2986/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2996 U$$2996/A U$$3000/B VGND VGND VPWR VPWR U$$2996/X sky130_fd_sc_hd__xor2_1
XANTENNA_290 _214_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_44_5 U$$2090/X U$$2223/X VGND VGND VPWR VPWR dadda_fa_2_45_4/A dadda_fa_3_44_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_970 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_50_4 U$$1703/X U$$1836/X U$$1969/X VGND VGND VPWR VPWR dadda_fa_2_51_1/CIN
+ dadda_fa_2_50_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$808 U$$808/A U$$810/B VGND VGND VPWR VPWR U$$808/X sky130_fd_sc_hd__xor2_1
XU$$819 U$$956/A1 U$$819/A2 U$$819/B1 U$$819/B2 VGND VGND VPWR VPWR U$$820/A sky130_fd_sc_hd__a22o_1
XFILLER_56_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_43_3 U$$1290/X U$$1423/X U$$1556/X VGND VGND VPWR VPWR dadda_fa_2_44_3/CIN
+ dadda_fa_2_43_5/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_20_2 dadda_fa_4_20_2/A dadda_fa_4_20_2/B dadda_ha_3_20_3/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_21_0/CIN dadda_fa_5_20_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_97_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_13_1 U$$432/X U$$565/X U$$698/X VGND VGND VPWR VPWR dadda_fa_5_14_0/B
+ dadda_fa_5_13_1/B sky130_fd_sc_hd__fa_1
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1708 _552_/Q VGND VGND VPWR VPWR U$$3157/B1 sky130_fd_sc_hd__buf_4
XFILLER_137_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_58_3 dadda_fa_3_58_3/A dadda_fa_3_58_3/B dadda_fa_3_58_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_1/B dadda_fa_4_58_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2204 U$$2478/A1 U$$2242/A2 U$$2343/A1 U$$2242/B2 VGND VGND VPWR VPWR U$$2205/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2215 U$$2215/A U$$2263/B VGND VGND VPWR VPWR U$$2215/X sky130_fd_sc_hd__xor2_1
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2226 U$$3320/B1 U$$2302/A2 U$$719/B1 U$$2302/B2 VGND VGND VPWR VPWR U$$2227/A
+ sky130_fd_sc_hd__a22o_1
XU$$2237 U$$2237/A U$$2243/B VGND VGND VPWR VPWR U$$2237/X sky130_fd_sc_hd__xor2_1
XU$$1503 U$$1503/A U$$1507/A VGND VGND VPWR VPWR U$$1503/X sky130_fd_sc_hd__xor2_1
XU$$2248 U$$4027/B1 U$$2248/A2 U$$3346/A1 U$$2248/B2 VGND VGND VPWR VPWR U$$2249/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2259 U$$2259/A U$$2269/B VGND VGND VPWR VPWR U$$2259/X sky130_fd_sc_hd__xor2_1
XU$$1514 U$$1514/A U$$1558/B VGND VGND VPWR VPWR U$$1514/X sky130_fd_sc_hd__xor2_1
XU$$1525 U$$840/A1 U$$1553/A2 U$$705/A1 U$$1553/B2 VGND VGND VPWR VPWR U$$1526/A sky130_fd_sc_hd__a22o_1
XFILLER_37_1104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1536 U$$1536/A U$$1578/B VGND VGND VPWR VPWR U$$1536/X sky130_fd_sc_hd__xor2_1
XFILLER_16_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1547 U$$451/A1 U$$1561/A2 U$$999/B1 U$$1561/B2 VGND VGND VPWR VPWR U$$1548/A sky130_fd_sc_hd__a22o_1
XFILLER_203_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1558 U$$1558/A U$$1558/B VGND VGND VPWR VPWR U$$1558/X sky130_fd_sc_hd__xor2_1
XFILLER_30_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1569 U$$1843/A1 U$$1577/A2 U$$749/A1 U$$1577/B2 VGND VGND VPWR VPWR U$$1570/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_228_ _353_/CLK _228_/D VGND VGND VPWR VPWR _228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_84_0_1856 VGND VGND VPWR VPWR dadda_fa_1_84_0/A dadda_fa_1_84_0_1856/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_97_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_3 dadda_fa_2_60_3/A dadda_fa_2_60_3/B dadda_fa_2_60_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/B dadda_fa_3_60_3/B sky130_fd_sc_hd__fa_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater403 U$$819/A2 VGND VGND VPWR VPWR U$$783/A2 sky130_fd_sc_hd__buf_4
Xrepeater414 U$$682/A2 VGND VGND VPWR VPWR U$$650/A2 sky130_fd_sc_hd__buf_4
XFILLER_211_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater425 U$$491/A2 VGND VGND VPWR VPWR U$$457/A2 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_2_53_2 dadda_fa_2_53_2/A dadda_fa_2_53_2/B dadda_fa_2_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/A dadda_fa_3_53_3/A sky130_fd_sc_hd__fa_1
Xrepeater436 U$$4196/A2 VGND VGND VPWR VPWR U$$4182/A2 sky130_fd_sc_hd__buf_4
XFILLER_84_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_832 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater447 U$$4065/A2 VGND VGND VPWR VPWR U$$4029/A2 sky130_fd_sc_hd__buf_6
XFILLER_38_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4140 U$$4140/A1 U$$4140/A2 U$$4140/B1 U$$4140/B2 VGND VGND VPWR VPWR U$$4141/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater458 U$$3840/X VGND VGND VPWR VPWR U$$3910/A2 sky130_fd_sc_hd__buf_6
XU$$4151 U$$4151/A U$$4183/B VGND VGND VPWR VPWR U$$4151/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1001 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_30_1 dadda_fa_5_30_1/A dadda_fa_5_30_1/B dadda_fa_5_30_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_31_0/B dadda_fa_7_30_0/A sky130_fd_sc_hd__fa_1
Xrepeater469 U$$3703/X VGND VGND VPWR VPWR U$$3805/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_46_1 U$$3158/X U$$3208/B input197/X VGND VGND VPWR VPWR dadda_fa_3_47_0/CIN
+ dadda_fa_3_46_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_93_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4162 _574_/Q U$$4174/A2 _575_/Q U$$4174/B2 VGND VGND VPWR VPWR U$$4163/A sky130_fd_sc_hd__a22o_1
XU$$4173 U$$4173/A U$$4175/B VGND VGND VPWR VPWR U$$4173/X sky130_fd_sc_hd__xor2_1
XU$$4184 U$$4184/A1 U$$4196/A2 U$$4186/A1 U$$4196/B2 VGND VGND VPWR VPWR U$$4185/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_23_0 dadda_fa_5_23_0/A dadda_fa_5_23_0/B dadda_fa_5_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_24_0/A dadda_fa_6_23_0/CIN sky130_fd_sc_hd__fa_2
XU$$4195 U$$4195/A U$$4197/B VGND VGND VPWR VPWR U$$4195/X sky130_fd_sc_hd__xor2_1
XFILLER_81_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3450 U$$3450/A U$$3498/B VGND VGND VPWR VPWR U$$3450/X sky130_fd_sc_hd__xor2_1
XFILLER_207_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3461 U$$3735/A1 U$$3559/A2 U$$3735/B1 U$$3559/B2 VGND VGND VPWR VPWR U$$3462/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_39_0 U$$1149/X U$$1282/X U$$1415/X VGND VGND VPWR VPWR dadda_fa_3_40_0/B
+ dadda_fa_3_39_2/B sky130_fd_sc_hd__fa_1
XU$$3472 U$$3472/A U$$3506/B VGND VGND VPWR VPWR U$$3472/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_334 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3483 _577_/Q U$$3519/A2 U$$3485/A1 U$$3519/B2 VGND VGND VPWR VPWR U$$3484/A sky130_fd_sc_hd__a22o_1
XFILLER_20_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3494 U$$3494/A U$$3498/B VGND VGND VPWR VPWR U$$3494/X sky130_fd_sc_hd__xor2_1
XU$$2760 U$$3717/B1 U$$2788/A2 _559_/Q U$$2788/B2 VGND VGND VPWR VPWR U$$2761/A sky130_fd_sc_hd__a22o_1
XFILLER_206_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2771 U$$2771/A U$$2827/B VGND VGND VPWR VPWR U$$2771/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2782 U$$3876/B1 U$$2788/A2 U$$3056/B1 U$$2788/B2 VGND VGND VPWR VPWR U$$2783/A
+ sky130_fd_sc_hd__a22o_1
XU$$2793 U$$2793/A U$$2795/B VGND VGND VPWR VPWR U$$2793/X sky130_fd_sc_hd__xor2_1
XFILLER_178_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1787_1725 VGND VGND VPWR VPWR U$$1787_1725/HI U$$1787/A1 sky130_fd_sc_hd__conb_1
XFILLER_179_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_68_2 dadda_fa_4_68_2/A dadda_fa_4_68_2/B dadda_fa_4_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/CIN dadda_fa_5_68_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput206 c[54] VGND VGND VPWR VPWR input206/X sky130_fd_sc_hd__clkbuf_4
Xinput217 c[64] VGND VGND VPWR VPWR input217/X sky130_fd_sc_hd__clkbuf_1
Xinput228 c[74] VGND VGND VPWR VPWR input228/X sky130_fd_sc_hd__clkbuf_4
XTAP_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1030 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput239 c[84] VGND VGND VPWR VPWR input239/X sky130_fd_sc_hd__clkbuf_2
Xfinal_adder.U$$700 final_adder.U$$700/A final_adder.U$$700/B VGND VGND VPWR VPWR
+ _246_/D sky130_fd_sc_hd__xor2_1
XTAP_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_38_0 dadda_fa_7_38_0/A dadda_fa_7_38_0/B dadda_fa_7_38_0/CIN VGND VGND
+ VPWR VPWR _463_/D _334_/D sky130_fd_sc_hd__fa_1
XFILLER_57_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$711 final_adder.U$$711/A final_adder.U$$711/B VGND VGND VPWR VPWR
+ _257_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$722 final_adder.U$$722/A final_adder.U$$722/B VGND VGND VPWR VPWR
+ _268_/D sky130_fd_sc_hd__xor2_1
XTAP_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$733 final_adder.U$$733/A final_adder.U$$733/B VGND VGND VPWR VPWR
+ _279_/D sky130_fd_sc_hd__xor2_4
XTAP_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$744 final_adder.U$$744/A final_adder.U$$744/B VGND VGND VPWR VPWR
+ _290_/D sky130_fd_sc_hd__xor2_4
XFILLER_5_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$605 U$$605/A U$$613/B VGND VGND VPWR VPWR U$$605/X sky130_fd_sc_hd__xor2_1
XFILLER_17_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater970 U$$3424/A VGND VGND VPWR VPWR U$$3369/B sky130_fd_sc_hd__buf_8
Xrepeater981 U$$3288/A VGND VGND VPWR VPWR U$$3286/B sky130_fd_sc_hd__buf_6
XFILLER_72_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$616 U$$68/A1 U$$616/A2 U$$70/A1 U$$616/B2 VGND VGND VPWR VPWR U$$617/A sky130_fd_sc_hd__a22o_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_41_0 U$$89/X U$$222/X U$$355/X VGND VGND VPWR VPWR dadda_fa_2_42_3/B dadda_fa_2_41_5/A
+ sky130_fd_sc_hd__fa_1
XU$$627 U$$627/A U$$627/B VGND VGND VPWR VPWR U$$627/X sky130_fd_sc_hd__xor2_1
XFILLER_99_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater992 _661_/Q VGND VGND VPWR VPWR U$$3145/B sky130_fd_sc_hd__buf_6
XFILLER_84_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$638 U$$912/A1 U$$650/A2 U$$912/B1 U$$650/B2 VGND VGND VPWR VPWR U$$639/A sky130_fd_sc_hd__a22o_1
XFILLER_112_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$649 U$$649/A U$$651/B VGND VGND VPWR VPWR U$$649/X sky130_fd_sc_hd__xor2_1
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2746_1740 VGND VGND VPWR VPWR U$$2746_1740/HI U$$2746/A1 sky130_fd_sc_hd__conb_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_20 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1001 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1072 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1505 U$$4442/A1 VGND VGND VPWR VPWR U$$4305/A1 sky130_fd_sc_hd__buf_4
Xrepeater1516 _575_/Q VGND VGND VPWR VPWR U$$4436/B1 sky130_fd_sc_hd__buf_6
XFILLER_137_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1527 U$$3475/B1 VGND VGND VPWR VPWR U$$463/A1 sky130_fd_sc_hd__buf_4
XFILLER_193_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1538 U$$4160/A1 VGND VGND VPWR VPWR U$$3475/A1 sky130_fd_sc_hd__buf_4
Xrepeater1549 U$$731/A1 VGND VGND VPWR VPWR U$$729/B1 sky130_fd_sc_hd__buf_4
XFILLER_158_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_70_2 dadda_fa_3_70_2/A dadda_fa_3_70_2/B dadda_fa_3_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_1/A dadda_fa_4_70_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_0_72_0_1851 VGND VGND VPWR VPWR dadda_fa_0_72_0/A dadda_fa_0_72_0_1851/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_63_1 dadda_fa_3_63_1/A dadda_fa_3_63_1/B dadda_fa_3_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_0/CIN dadda_fa_4_63_2/A sky130_fd_sc_hd__fa_1
XFILLER_94_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_40_0 dadda_fa_6_40_0/A dadda_fa_6_40_0/B dadda_fa_6_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_41_0/B dadda_fa_7_40_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_56_0 dadda_fa_3_56_0/A dadda_fa_3_56_0/B dadda_fa_3_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_0/B dadda_fa_4_56_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2001 U$$2001/A U$$2003/B VGND VGND VPWR VPWR U$$2001/X sky130_fd_sc_hd__xor2_1
XU$$2012 U$$368/A1 U$$2028/A2 U$$96/A1 U$$2028/B2 VGND VGND VPWR VPWR U$$2013/A sky130_fd_sc_hd__a22o_1
XFILLER_207_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2023 U$$2023/A U$$2029/B VGND VGND VPWR VPWR U$$2023/X sky130_fd_sc_hd__xor2_1
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2034 U$$2171/A1 U$$2038/A2 U$$392/A1 U$$2038/B2 VGND VGND VPWR VPWR U$$2035/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2045 U$$2045/A U$$2054/A VGND VGND VPWR VPWR U$$2045/X sky130_fd_sc_hd__xor2_1
XU$$1300 U$$1300/A U$$1310/B VGND VGND VPWR VPWR U$$1300/X sky130_fd_sc_hd__xor2_1
XU$$1311 U$$78/A1 U$$1355/A2 U$$2957/A1 U$$1355/B2 VGND VGND VPWR VPWR U$$1312/A sky130_fd_sc_hd__a22o_1
XU$$2056 _646_/Q VGND VGND VPWR VPWR U$$2058/B sky130_fd_sc_hd__inv_1
XU$$1322 U$$1322/A U$$1356/B VGND VGND VPWR VPWR U$$1322/X sky130_fd_sc_hd__xor2_1
XU$$2067 U$$2478/A1 U$$2115/A2 U$$2343/A1 U$$2115/B2 VGND VGND VPWR VPWR U$$2068/A
+ sky130_fd_sc_hd__a22o_1
XU$$2078 U$$2078/A U$$2110/B VGND VGND VPWR VPWR U$$2078/X sky130_fd_sc_hd__xor2_1
XU$$1333 U$$2838/B1 U$$1237/X U$$2705/A1 U$$1238/X VGND VGND VPWR VPWR U$$1334/A sky130_fd_sc_hd__a22o_1
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2089 U$$3320/B1 U$$2129/A2 U$$856/B1 U$$2129/B2 VGND VGND VPWR VPWR U$$2090/A
+ sky130_fd_sc_hd__a22o_1
XU$$1344 U$$1344/A U$$1369/A VGND VGND VPWR VPWR U$$1344/X sky130_fd_sc_hd__xor2_1
XU$$1355 U$$2725/A1 U$$1355/A2 U$$2588/B1 U$$1355/B2 VGND VGND VPWR VPWR U$$1356/A
+ sky130_fd_sc_hd__a22o_1
XU$$1366 U$$1366/A U$$1368/B VGND VGND VPWR VPWR U$$1366/X sky130_fd_sc_hd__xor2_1
XFILLER_149_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1377 U$$1377/A U$$1429/B VGND VGND VPWR VPWR U$$1377/X sky130_fd_sc_hd__xor2_1
XU$$1388 U$$2756/B1 U$$1424/A2 U$$840/B1 U$$1424/B2 VGND VGND VPWR VPWR U$$1389/A
+ sky130_fd_sc_hd__a22o_1
XU$$1399 U$$1399/A U$$1425/B VGND VGND VPWR VPWR U$$1399/X sky130_fd_sc_hd__xor2_1
XFILLER_176_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_113_0 dadda_fa_7_113_0/A dadda_fa_7_113_0/B dadda_fa_7_113_0/CIN VGND
+ VGND VPWR VPWR _538_/D _409_/D sky130_fd_sc_hd__fa_1
XFILLER_50_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_450 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_78_1 dadda_fa_5_78_1/A dadda_fa_5_78_1/B dadda_fa_5_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_79_0/B dadda_fa_7_78_0/A sky130_fd_sc_hd__fa_1
XFILLER_87_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$40 _464_/Q _336_/Q VGND VGND VPWR VPWR final_adder.U$$535/B1 final_adder.U$$662/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$51 _475_/Q _347_/Q VGND VGND VPWR VPWR final_adder.U$$179/B1 final_adder.U$$673/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3280 U$$3280/A U$$3288/A VGND VGND VPWR VPWR U$$3280/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$62 _486_/Q _358_/Q VGND VGND VPWR VPWR final_adder.U$$557/B1 final_adder.U$$684/A
+ sky130_fd_sc_hd__ha_1
XU$$3291 U$$3423/B U$$3291/B VGND VGND VPWR VPWR U$$3291/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$73 _497_/Q _369_/Q VGND VGND VPWR VPWR final_adder.U$$201/B1 final_adder.U$$695/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$84 _508_/Q _380_/Q VGND VGND VPWR VPWR final_adder.U$$579/B1 final_adder.U$$706/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$95 _519_/Q _391_/Q VGND VGND VPWR VPWR final_adder.U$$223/B1 final_adder.U$$717/A
+ sky130_fd_sc_hd__ha_1
XFILLER_34_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2590 _610_/Q U$$2600/A2 _611_/Q U$$2600/B2 VGND VGND VPWR VPWR U$$2591/A sky130_fd_sc_hd__a22o_1
XFILLER_22_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_80_1 dadda_fa_4_80_1/A dadda_fa_4_80_1/B dadda_fa_4_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/B dadda_fa_5_80_1/B sky130_fd_sc_hd__fa_1
XFILLER_119_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2737_1739 VGND VGND VPWR VPWR U$$2737_1739/HI U$$2737/B1 sky130_fd_sc_hd__conb_1
XFILLER_123_818 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_784 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_73_0 dadda_fa_4_73_0/A dadda_fa_4_73_0/B dadda_fa_4_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/A dadda_fa_5_73_1/A sky130_fd_sc_hd__fa_1
XFILLER_116_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_89_0 U$$1780/Y U$$1914/X U$$2047/X VGND VGND VPWR VPWR dadda_fa_2_90_3/CIN
+ dadda_fa_2_89_5/A sky130_fd_sc_hd__fa_1
XFILLER_135_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_927 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$541 final_adder.U$$668/A final_adder.U$$668/B final_adder.U$$541/B1
+ VGND VGND VPWR VPWR final_adder.U$$669/B sky130_fd_sc_hd__a21o_1
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_631_ _633_/CLK _631_/D VGND VGND VPWR VPWR _631_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$402 U$$676/A1 U$$408/A2 U$$676/B1 U$$408/B2 VGND VGND VPWR VPWR U$$403/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$563 final_adder.U$$690/A final_adder.U$$690/B final_adder.U$$563/B1
+ VGND VGND VPWR VPWR final_adder.U$$691/B sky130_fd_sc_hd__a21o_1
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$413 _623_/Q VGND VGND VPWR VPWR U$$413/Y sky130_fd_sc_hd__inv_1
XFILLER_205_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$424 U$$424/A U$$452/B VGND VGND VPWR VPWR U$$424/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$585 final_adder.U$$712/A final_adder.U$$712/B final_adder.U$$585/B1
+ VGND VGND VPWR VPWR final_adder.U$$713/B sky130_fd_sc_hd__a21o_1
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$435 U$$435/A1 U$$491/A2 U$$435/B1 U$$491/B2 VGND VGND VPWR VPWR U$$436/A sky130_fd_sc_hd__a22o_1
X_562_ _569_/CLK _562_/D VGND VGND VPWR VPWR _562_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$446 U$$446/A U$$452/B VGND VGND VPWR VPWR U$$446/X sky130_fd_sc_hd__xor2_1
XFILLER_45_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$457 U$$729/B1 U$$457/A2 U$$733/A1 U$$457/B2 VGND VGND VPWR VPWR U$$458/A sky130_fd_sc_hd__a22o_1
XU$$468 U$$468/A U$$500/B VGND VGND VPWR VPWR U$$468/X sky130_fd_sc_hd__xor2_1
XU$$479 U$$614/B1 U$$483/A2 U$$70/A1 U$$483/B2 VGND VGND VPWR VPWR U$$480/A sky130_fd_sc_hd__a22o_1
XFILLER_38_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_493_ _634_/CLK _493_/D VGND VGND VPWR VPWR _493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_450 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1302 U$$4218/A1 VGND VGND VPWR VPWR U$$4490/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_6_88_0 dadda_fa_6_88_0/A dadda_fa_6_88_0/B dadda_fa_6_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_89_0/B dadda_fa_7_88_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_931 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1313 _601_/Q VGND VGND VPWR VPWR U$$3805/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_78_0 dadda_ha_0_78_0/A U$$1094/X VGND VGND VPWR VPWR dadda_fa_2_79_0/A
+ dadda_fa_2_78_0/A sky130_fd_sc_hd__ha_1
Xrepeater1324 U$$785/B1 VGND VGND VPWR VPWR U$$648/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_5_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1335 U$$4484/A1 VGND VGND VPWR VPWR U$$2838/B1 sky130_fd_sc_hd__buf_4
Xrepeater1346 _597_/Q VGND VGND VPWR VPWR U$$4206/B1 sky130_fd_sc_hd__buf_6
XFILLER_4_441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1357 U$$368/A1 VGND VGND VPWR VPWR U$$94/A1 sky130_fd_sc_hd__buf_4
XFILLER_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1368 U$$4476/A1 VGND VGND VPWR VPWR U$$92/A1 sky130_fd_sc_hd__buf_4
Xrepeater1379 U$$4061/A1 VGND VGND VPWR VPWR U$$910/A1 sky130_fd_sc_hd__buf_4
XFILLER_180_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_835 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1029 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_985 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$980 U$$980/A U$$980/B VGND VGND VPWR VPWR U$$980/X sky130_fd_sc_hd__xor2_1
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$991 U$$991/A1 U$$995/A2 U$$34/A1 U$$995/B2 VGND VGND VPWR VPWR U$$992/A sky130_fd_sc_hd__a22o_1
XU$$1130 U$$993/A1 U$$1190/A2 U$$856/B1 U$$1190/B2 VGND VGND VPWR VPWR U$$1131/A sky130_fd_sc_hd__a22o_1
XFILLER_91_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1141 U$$1141/A U$$1147/B VGND VGND VPWR VPWR U$$1141/X sky130_fd_sc_hd__xor2_1
XU$$1152 U$$330/A1 U$$1194/A2 U$$58/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1153/A sky130_fd_sc_hd__a22o_1
XU$$1163 U$$1163/A U$$1191/B VGND VGND VPWR VPWR U$$1163/X sky130_fd_sc_hd__xor2_1
XU$$1174 U$$78/A1 U$$1176/A2 U$$80/A1 U$$1176/B2 VGND VGND VPWR VPWR U$$1175/A sky130_fd_sc_hd__a22o_1
XFILLER_149_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1185 U$$1185/A U$$1225/B VGND VGND VPWR VPWR U$$1185/X sky130_fd_sc_hd__xor2_1
XFILLER_188_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1196 U$$2838/B1 U$$1208/A2 U$$2705/A1 U$$1208/B2 VGND VGND VPWR VPWR U$$1197/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_90_0 dadda_fa_5_90_0/A dadda_fa_5_90_0/B dadda_fa_5_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_91_0/A dadda_fa_6_90_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_75_6 U$$4014/X U$$4147/X U$$4280/X VGND VGND VPWR VPWR dadda_fa_2_76_2/B
+ dadda_fa_2_75_5/B sky130_fd_sc_hd__fa_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_5 input221/X dadda_fa_1_68_5/B dadda_fa_1_68_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_69_2/A dadda_fa_2_68_5/A sky130_fd_sc_hd__fa_2
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_108 _179_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_119 _289_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2600_1736 VGND VGND VPWR VPWR U$$2600_1736/HI U$$2600/B1 sky130_fd_sc_hd__conb_1
XFILLER_120_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_120_0 dadda_fa_6_120_0/A dadda_fa_6_120_0/B dadda_fa_6_120_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_121_0/B dadda_fa_7_120_0/CIN sky130_fd_sc_hd__fa_1
XTAP_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_4 U$$1729/X U$$1862/X U$$1995/X VGND VGND VPWR VPWR dadda_fa_1_64_6/CIN
+ dadda_fa_1_63_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_40_3 dadda_fa_3_40_3/A dadda_fa_3_40_3/B dadda_fa_3_40_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_1/B dadda_fa_4_40_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$360 final_adder.U$$360/A final_adder.U$$360/B VGND VGND VPWR VPWR
+ final_adder.U$$372/B sky130_fd_sc_hd__and2_1
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$371 final_adder.U$$370/A final_adder.U$$357/X final_adder.U$$359/X
+ VGND VGND VPWR VPWR final_adder.U$$371/X sky130_fd_sc_hd__a21o_1
XU$$210 U$$210/A U$$216/B VGND VGND VPWR VPWR U$$210/X sky130_fd_sc_hd__xor2_1
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_614_ _615_/CLK _614_/D VGND VGND VPWR VPWR _614_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_33_2 dadda_fa_3_33_2/A dadda_fa_3_33_2/B dadda_fa_3_33_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_1/A dadda_fa_4_33_2/B sky130_fd_sc_hd__fa_1
XU$$221 U$$358/A1 U$$263/A2 U$$86/A1 U$$263/B2 VGND VGND VPWR VPWR U$$222/A sky130_fd_sc_hd__a22o_1
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$393 final_adder.U$$356/B final_adder.U$$654/B final_adder.U$$329/X
+ VGND VGND VPWR VPWR final_adder.U$$662/B sky130_fd_sc_hd__a21o_2
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$232 U$$232/A U$$232/B VGND VGND VPWR VPWR U$$232/X sky130_fd_sc_hd__xor2_1
XU$$243 U$$515/B1 U$$249/A2 U$$517/B1 U$$249/B2 VGND VGND VPWR VPWR U$$244/A sky130_fd_sc_hd__a22o_1
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$254 U$$254/A U$$264/B VGND VGND VPWR VPWR U$$254/X sky130_fd_sc_hd__xor2_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$265 U$$676/A1 U$$141/X U$$676/B1 U$$142/X VGND VGND VPWR VPWR U$$266/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_26_1 U$$1522/X U$$1655/X U$$1788/X VGND VGND VPWR VPWR dadda_fa_4_27_0/CIN
+ dadda_fa_4_26_2/A sky130_fd_sc_hd__fa_1
XFILLER_72_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_545_ _547_/CLK _545_/D VGND VGND VPWR VPWR _545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$276 _621_/Q VGND VGND VPWR VPWR U$$276/Y sky130_fd_sc_hd__inv_1
XU$$287 U$$287/A U$$319/B VGND VGND VPWR VPWR U$$287/X sky130_fd_sc_hd__xor2_1
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$298 U$$22/B1 U$$308/A2 U$$26/A1 U$$308/B2 VGND VGND VPWR VPWR U$$299/A sky130_fd_sc_hd__a22o_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_19_0 U$$45/X U$$178/X U$$311/X VGND VGND VPWR VPWR dadda_fa_4_20_0/CIN
+ dadda_fa_4_19_2/A sky130_fd_sc_hd__fa_1
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_476_ _476_/CLK _476_/D VGND VGND VPWR VPWR _476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4 U$$2/Y U$$1/A U$$4/A3 U$$3/X U$$0/Y VGND VGND VPWR VPWR U$$4/X sky130_fd_sc_hd__a32o_4
XFILLER_51_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1110 _635_/Q VGND VGND VPWR VPWR U$$1370/A sky130_fd_sc_hd__buf_4
Xrepeater1121 U$$1078/B VGND VGND VPWR VPWR U$$996/B sky130_fd_sc_hd__buf_6
Xoutput307 _170_/Q VGND VGND VPWR VPWR o[2] sky130_fd_sc_hd__buf_2
Xoutput318 _171_/Q VGND VGND VPWR VPWR o[3] sky130_fd_sc_hd__buf_2
XFILLER_126_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1132 U$$897/B VGND VGND VPWR VPWR U$$907/B sky130_fd_sc_hd__buf_6
Xoutput329 _172_/Q VGND VGND VPWR VPWR o[4] sky130_fd_sc_hd__buf_2
XFILLER_141_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1143 U$$821/A VGND VGND VPWR VPWR U$$816/B sky130_fd_sc_hd__buf_8
XFILLER_142_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1154 U$$685/A VGND VGND VPWR VPWR U$$669/B sky130_fd_sc_hd__buf_6
XFILLER_142_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1165 U$$335/B VGND VGND VPWR VPWR U$$309/B sky130_fd_sc_hd__buf_6
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_85_5 dadda_fa_2_85_5/A dadda_fa_2_85_5/B dadda_fa_2_85_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_2/A dadda_fa_4_85_0/A sky130_fd_sc_hd__fa_2
Xrepeater1176 U$$216/B VGND VGND VPWR VPWR U$$180/B sky130_fd_sc_hd__clkbuf_8
XFILLER_99_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1187 U$$117/B VGND VGND VPWR VPWR U$$85/B sky130_fd_sc_hd__buf_6
Xrepeater1198 _615_/Q VGND VGND VPWR VPWR U$$2872/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_78_4 dadda_fa_2_78_4/A dadda_fa_2_78_4/B dadda_fa_2_78_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/CIN dadda_fa_3_78_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_101_3 U$$3800/X U$$3933/X U$$4066/X VGND VGND VPWR VPWR dadda_fa_3_102_2/CIN
+ dadda_fa_4_101_0/A sky130_fd_sc_hd__fa_1
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_115_1 dadda_fa_5_115_1/A dadda_fa_5_115_1/B dadda_fa_5_115_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_116_0/B dadda_fa_7_115_0/A sky130_fd_sc_hd__fa_1
XFILLER_117_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_108_0 dadda_fa_5_108_0/A dadda_fa_5_108_0/B dadda_fa_5_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_109_0/A dadda_fa_6_108_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_80_4 U$$2694/X U$$2827/X U$$2960/X VGND VGND VPWR VPWR dadda_fa_2_81_2/A
+ dadda_fa_2_80_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_73_3 U$$3079/X U$$3212/X U$$3345/X VGND VGND VPWR VPWR dadda_fa_2_74_1/B
+ dadda_fa_2_73_4/B sky130_fd_sc_hd__fa_1
XFILLER_154_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_50_2 dadda_fa_4_50_2/A dadda_fa_4_50_2/B dadda_fa_4_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/CIN dadda_fa_5_50_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_24_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_66_2 U$$3331/X U$$3464/X U$$3597/X VGND VGND VPWR VPWR dadda_fa_2_67_1/A
+ dadda_fa_2_66_4/A sky130_fd_sc_hd__fa_1
XFILLER_115_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4413_1785 VGND VGND VPWR VPWR U$$4413_1785/HI U$$4413/B sky130_fd_sc_hd__conb_1
XFILLER_86_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_43_1 dadda_fa_4_43_1/A dadda_fa_4_43_1/B dadda_fa_4_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/B dadda_fa_5_43_1/B sky130_fd_sc_hd__fa_1
XFILLER_46_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_59_1 U$$1987/X U$$2120/X U$$2253/X VGND VGND VPWR VPWR dadda_fa_2_60_0/CIN
+ dadda_fa_2_59_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_20_0 dadda_fa_7_20_0/A dadda_fa_7_20_0/B dadda_fa_7_20_0/CIN VGND VGND
+ VPWR VPWR _445_/D _316_/D sky130_fd_sc_hd__fa_1
XFILLER_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_36_0 dadda_fa_4_36_0/A dadda_fa_4_36_0/B dadda_fa_4_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/A dadda_fa_5_36_1/A sky130_fd_sc_hd__fa_1
XFILLER_6_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1092 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_330_ _458_/CLK _330_/D VGND VGND VPWR VPWR _330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_955 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _519_/CLK _261_/D VGND VGND VPWR VPWR _261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_192_ _207_/CLK _192_/D VGND VGND VPWR VPWR _192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_20 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_75 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1513_1721 VGND VGND VPWR VPWR U$$1513_1721/HI U$$1513/A1 sky130_fd_sc_hd__conb_1
XFILLER_159_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_88_3 dadda_fa_3_88_3/A dadda_fa_3_88_3/B dadda_fa_3_88_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_1/B dadda_fa_4_88_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_97_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4503 U$$4503/A U$$4503/B VGND VGND VPWR VPWR U$$4503/X sky130_fd_sc_hd__xor2_1
XU$$4514 U$$4514/A1 U$$4388/X U$$4516/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4515/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_61_1 U$$528/X U$$661/X U$$794/X VGND VGND VPWR VPWR dadda_fa_1_62_6/A
+ dadda_fa_1_61_8/A sky130_fd_sc_hd__fa_1
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$17 U$$17/A U$$9/B VGND VGND VPWR VPWR U$$17/X sky130_fd_sc_hd__xor2_1
XU$$3802 U$$3802/A U$$3804/B VGND VGND VPWR VPWR U$$3802/X sky130_fd_sc_hd__xor2_1
XU$$3813 U$$4087/A1 U$$3703/X U$$4087/B1 U$$3704/X VGND VGND VPWR VPWR U$$3814/A sky130_fd_sc_hd__a22o_1
XU$$28 U$$28/A1 U$$52/A2 U$$30/A1 U$$52/B2 VGND VGND VPWR VPWR U$$29/A sky130_fd_sc_hd__a22o_1
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_54_0 U$$115/X U$$248/X U$$381/X VGND VGND VPWR VPWR dadda_fa_1_55_8/A
+ dadda_fa_1_54_8/CIN sky130_fd_sc_hd__fa_1
XU$$3824 U$$3824/A U$$3832/B VGND VGND VPWR VPWR U$$3824/X sky130_fd_sc_hd__xor2_1
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3835 U$$3835/A VGND VGND VPWR VPWR U$$3835/Y sky130_fd_sc_hd__inv_1
XU$$39 U$$39/A U$$3/A VGND VGND VPWR VPWR U$$39/X sky130_fd_sc_hd__xor2_1
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3846 U$$4394/A1 U$$3910/A2 _554_/Q U$$3910/B2 VGND VGND VPWR VPWR U$$3847/A sky130_fd_sc_hd__a22o_1
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$190 final_adder.U$$685/A final_adder.U$$684/A VGND VGND VPWR VPWR
+ final_adder.U$$286/A sky130_fd_sc_hd__and2_1
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3857 U$$3857/A U$$3965/B VGND VGND VPWR VPWR U$$3857/X sky130_fd_sc_hd__xor2_1
XU$$3868 _564_/Q U$$3958/A2 _565_/Q U$$3958/B2 VGND VGND VPWR VPWR U$$3869/A sky130_fd_sc_hd__a22o_1
XU$$3879 U$$3879/A U$$3917/B VGND VGND VPWR VPWR U$$3879/X sky130_fd_sc_hd__xor2_1
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_777 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_528_ _566_/CLK _528_/D VGND VGND VPWR VPWR _528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_19 _281_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_459_ _463_/CLK _459_/D VGND VGND VPWR VPWR _459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_90_3 U$$4443/X input246/X dadda_fa_2_90_3/CIN VGND VGND VPWR VPWR dadda_fa_3_91_1/B
+ dadda_fa_3_90_3/B sky130_fd_sc_hd__fa_1
XFILLER_126_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_120_0_1871 VGND VGND VPWR VPWR dadda_fa_4_120_0/A dadda_fa_4_120_0_1871/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_83_2 dadda_fa_2_83_2/A dadda_fa_2_83_2/B dadda_fa_2_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/A dadda_fa_3_83_3/A sky130_fd_sc_hd__fa_1
XFILLER_138_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_60_1 dadda_fa_5_60_1/A dadda_fa_5_60_1/B dadda_fa_5_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_61_0/B dadda_fa_7_60_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_76_1 dadda_fa_2_76_1/A dadda_fa_2_76_1/B dadda_fa_2_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_0/CIN dadda_fa_3_76_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_53_0 dadda_fa_5_53_0/A dadda_fa_5_53_0/B dadda_fa_5_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_54_0/A dadda_fa_6_53_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_141_297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_69_0 dadda_fa_2_69_0/A dadda_fa_2_69_0/B dadda_fa_2_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_0/B dadda_fa_3_69_2/B sky130_fd_sc_hd__fa_1
XFILLER_29_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_52_8 U$$3569/X U$$3613/B input204/X VGND VGND VPWR VPWR dadda_fa_2_53_3/A
+ dadda_fa_3_52_0/A sky130_fd_sc_hd__fa_1
XFILLER_3_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_98_2 dadda_fa_4_98_2/A dadda_fa_4_98_2/B dadda_fa_4_98_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/CIN dadda_fa_5_98_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_164_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_68_0 dadda_fa_7_68_0/A dadda_fa_7_68_0/B dadda_fa_7_68_0/CIN VGND VGND
+ VPWR VPWR _493_/D _364_/D sky130_fd_sc_hd__fa_1
XFILLER_79_808 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_71_0 U$$2144/X U$$2277/X U$$2410/X VGND VGND VPWR VPWR dadda_fa_2_72_0/B
+ dadda_fa_2_71_3/B sky130_fd_sc_hd__fa_1
XFILLER_143_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3109 U$$3109/A U$$3111/B VGND VGND VPWR VPWR U$$3109/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2408 U$$2408/A U$$2442/B VGND VGND VPWR VPWR U$$2408/X sky130_fd_sc_hd__xor2_1
XU$$2419 U$$3652/A1 U$$2423/A2 U$$914/A1 U$$2423/B2 VGND VGND VPWR VPWR U$$2420/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1707 U$$1707/A U$$1711/B VGND VGND VPWR VPWR U$$1707/X sky130_fd_sc_hd__xor2_1
XFILLER_27_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1718 U$$896/A1 U$$1718/A2 U$$896/B1 U$$1718/B2 VGND VGND VPWR VPWR U$$1719/A sky130_fd_sc_hd__a22o_1
XU$$1729 U$$1729/A U$$1737/B VGND VGND VPWR VPWR U$$1729/X sky130_fd_sc_hd__xor2_1
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_616 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_313_ _441_/CLK _313_/D VGND VGND VPWR VPWR _313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_244_ _372_/CLK _244_/D VGND VGND VPWR VPWR _244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput17 a[24] VGND VGND VPWR VPWR _640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput28 a[34] VGND VGND VPWR VPWR _650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput39 a[44] VGND VGND VPWR VPWR _660_/D sky130_fd_sc_hd__clkbuf_1
X_175_ _428_/CLK _175_/D VGND VGND VPWR VPWR _175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_93_1 dadda_fa_3_93_1/A dadda_fa_3_93_1/B dadda_fa_3_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_0/CIN dadda_fa_4_93_2/A sky130_fd_sc_hd__fa_1
XFILLER_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_70_0 dadda_fa_6_70_0/A dadda_fa_6_70_0/B dadda_fa_6_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_71_0/B dadda_fa_7_70_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_86_0 dadda_fa_3_86_0/A dadda_fa_3_86_0/B dadda_fa_3_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_0/B dadda_fa_4_86_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_184_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater607 U$$1511/X VGND VGND VPWR VPWR U$$1607/A2 sky130_fd_sc_hd__buf_4
XFILLER_81_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater618 U$$1478/A2 VGND VGND VPWR VPWR U$$1442/A2 sky130_fd_sc_hd__buf_4
XU$$4300 U$$4300/A U$$4348/B VGND VGND VPWR VPWR U$$4300/X sky130_fd_sc_hd__xor2_1
XFILLER_38_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater629 U$$1367/A2 VGND VGND VPWR VPWR U$$1355/A2 sky130_fd_sc_hd__buf_6
XFILLER_65_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4311 U$$4446/B1 U$$4311/A2 U$$4450/A1 U$$4311/B2 VGND VGND VPWR VPWR U$$4312/A
+ sky130_fd_sc_hd__a22o_1
XU$$4322 U$$4322/A U$$4322/B VGND VGND VPWR VPWR U$$4322/X sky130_fd_sc_hd__xor2_1
XFILLER_77_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4333 U$$4470/A1 U$$4335/A2 U$$4333/B1 U$$4333/B2 VGND VGND VPWR VPWR U$$4334/A
+ sky130_fd_sc_hd__a22o_1
XU$$4344 U$$4344/A U$$4350/B VGND VGND VPWR VPWR U$$4344/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4355 U$$4490/B1 U$$4369/A2 U$$4355/B1 U$$4369/B2 VGND VGND VPWR VPWR U$$4356/A
+ sky130_fd_sc_hd__a22o_1
XU$$3610 U$$4158/A1 U$$3612/A2 U$$4160/A1 U$$3612/B2 VGND VGND VPWR VPWR U$$3611/A
+ sky130_fd_sc_hd__a22o_1
XU$$3621 U$$3621/A U$$3663/B VGND VGND VPWR VPWR U$$3621/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_48_5 dadda_fa_2_48_5/A dadda_fa_2_48_5/B dadda_fa_2_48_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_2/A dadda_fa_4_48_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_115_0 U$$3961/X U$$4094/X U$$4227/X VGND VGND VPWR VPWR dadda_fa_5_116_0/A
+ dadda_fa_5_115_1/A sky130_fd_sc_hd__fa_1
XU$$4366 U$$4366/A U$$4384/A VGND VGND VPWR VPWR U$$4366/X sky130_fd_sc_hd__xor2_1
XFILLER_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4377 U$$4514/A1 U$$4381/A2 U$$4516/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4378/A
+ sky130_fd_sc_hd__a22o_1
XU$$3632 U$$3769/A1 U$$3696/A2 U$$3769/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3633/A
+ sky130_fd_sc_hd__a22o_1
XU$$4388 U$$4386/Y U$$4388/A2 U$$4384/A U$$4387/X U$$4384/Y VGND VGND VPWR VPWR U$$4388/X
+ sky130_fd_sc_hd__a32o_1
XU$$3643 U$$3643/A U$$3675/B VGND VGND VPWR VPWR U$$3643/X sky130_fd_sc_hd__xor2_1
XFILLER_203_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3654 U$$3789/B1 U$$3664/A2 U$$3791/B1 U$$3664/B2 VGND VGND VPWR VPWR U$$3655/A
+ sky130_fd_sc_hd__a22o_1
XU$$4399 U$$4399/A U$$4399/B VGND VGND VPWR VPWR U$$4399/X sky130_fd_sc_hd__xor2_1
XU$$3665 U$$3665/A U$$3671/B VGND VGND VPWR VPWR U$$3665/X sky130_fd_sc_hd__xor2_1
XFILLER_19_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2920 U$$2920/A U$$2944/B VGND VGND VPWR VPWR U$$2920/X sky130_fd_sc_hd__xor2_1
XU$$2931 U$$4436/B1 U$$2973/A2 U$$4301/B1 U$$2973/B2 VGND VGND VPWR VPWR U$$2932/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_387 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3676 U$$4087/A1 U$$3688/A2 U$$4087/B1 U$$3688/B2 VGND VGND VPWR VPWR U$$3677/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3687 U$$3687/A U$$3699/A VGND VGND VPWR VPWR U$$3687/X sky130_fd_sc_hd__xor2_1
XFILLER_18_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2942 U$$2942/A U$$2944/B VGND VGND VPWR VPWR U$$2942/X sky130_fd_sc_hd__xor2_1
XU$$2953 U$$4186/A1 U$$2959/A2 U$$4051/A1 U$$2959/B2 VGND VGND VPWR VPWR U$$2954/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_495 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3698 U$$3698/A VGND VGND VPWR VPWR U$$3698/Y sky130_fd_sc_hd__inv_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2964 U$$2964/A U$$2966/B VGND VGND VPWR VPWR U$$2964/X sky130_fd_sc_hd__xor2_1
XU$$2975 U$$4482/A1 U$$2881/X U$$4208/B1 U$$2882/X VGND VGND VPWR VPWR U$$2976/A sky130_fd_sc_hd__a22o_1
XU$$2986 U$$2986/A U$$2988/B VGND VGND VPWR VPWR U$$2986/X sky130_fd_sc_hd__xor2_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2997 U$$3269/B1 U$$2997/A2 _609_/Q U$$2997/B2 VGND VGND VPWR VPWR U$$2998/A sky130_fd_sc_hd__a22o_1
XFILLER_33_465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_291 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_999 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_982 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_50_5 U$$2102/X U$$2235/X U$$2368/X VGND VGND VPWR VPWR dadda_fa_2_51_2/A
+ dadda_fa_2_50_5/A sky130_fd_sc_hd__fa_1
XFILLER_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$809 U$$946/A1 U$$809/A2 U$$811/A1 U$$809/B2 VGND VGND VPWR VPWR U$$810/A sky130_fd_sc_hd__a22o_1
XFILLER_113_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3833_1756 VGND VGND VPWR VPWR U$$3833_1756/HI U$$3833/B1 sky130_fd_sc_hd__conb_1
XFILLER_58_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1709 _552_/Q VGND VGND VPWR VPWR U$$3844/A1 sky130_fd_sc_hd__buf_6
XFILLER_152_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2205 U$$2205/A U$$2241/B VGND VGND VPWR VPWR U$$2205/X sky130_fd_sc_hd__xor2_1
XFILLER_74_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2216 U$$435/A1 U$$2262/A2 U$$435/B1 U$$2262/B2 VGND VGND VPWR VPWR U$$2217/A sky130_fd_sc_hd__a22o_1
XFILLER_170_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2227 U$$2227/A U$$2303/B VGND VGND VPWR VPWR U$$2227/X sky130_fd_sc_hd__xor2_1
XU$$2238 U$$2375/A1 U$$2242/A2 U$$2375/B1 U$$2242/B2 VGND VGND VPWR VPWR U$$2239/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1504 U$$545/A1 U$$1374/X U$$1504/B1 U$$1375/X VGND VGND VPWR VPWR U$$1505/A sky130_fd_sc_hd__a22o_1
XU$$2249 U$$2249/A U$$2303/B VGND VGND VPWR VPWR U$$2249/X sky130_fd_sc_hd__xor2_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1515 U$$2746/B1 U$$1557/A2 U$$695/A1 U$$1557/B2 VGND VGND VPWR VPWR U$$1516/A
+ sky130_fd_sc_hd__a22o_1
XU$$1526 U$$1526/A U$$1554/B VGND VGND VPWR VPWR U$$1526/X sky130_fd_sc_hd__xor2_1
XFILLER_188_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1537 U$$3042/B1 U$$1577/A2 U$$2909/A1 U$$1577/B2 VGND VGND VPWR VPWR U$$1538/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1548 U$$1548/A U$$1562/B VGND VGND VPWR VPWR U$$1548/X sky130_fd_sc_hd__xor2_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1559 U$$600/A1 U$$1597/A2 U$$54/A1 U$$1597/B2 VGND VGND VPWR VPWR U$$1560/A sky130_fd_sc_hd__a22o_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_227_ _353_/CLK _227_/D VGND VGND VPWR VPWR _227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_4 dadda_fa_2_60_4/A dadda_fa_2_60_4/B dadda_fa_2_60_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/CIN dadda_fa_3_60_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater404 U$$809/A2 VGND VGND VPWR VPWR U$$819/A2 sky130_fd_sc_hd__buf_8
XFILLER_112_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater415 U$$552/X VGND VGND VPWR VPWR U$$682/A2 sky130_fd_sc_hd__buf_6
XFILLER_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater426 U$$499/A2 VGND VGND VPWR VPWR U$$483/A2 sky130_fd_sc_hd__buf_4
XFILLER_211_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_53_3 dadda_fa_2_53_3/A dadda_fa_2_53_3/B dadda_fa_2_53_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/B dadda_fa_3_53_3/B sky130_fd_sc_hd__fa_2
Xrepeater437 U$$4202/A2 VGND VGND VPWR VPWR U$$4196/A2 sky130_fd_sc_hd__buf_4
XFILLER_65_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater448 U$$4071/A2 VGND VGND VPWR VPWR U$$4065/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater459 U$$3958/A2 VGND VGND VPWR VPWR U$$3970/A2 sky130_fd_sc_hd__buf_4
XU$$4130 _558_/Q U$$4226/A2 U$$4269/A1 U$$4226/B2 VGND VGND VPWR VPWR U$$4131/A sky130_fd_sc_hd__a22o_1
XFILLER_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4141 U$$4141/A U$$4141/B VGND VGND VPWR VPWR U$$4141/X sky130_fd_sc_hd__xor2_1
XU$$4152 _569_/Q U$$4182/A2 U$$4154/A1 U$$4182/B2 VGND VGND VPWR VPWR U$$4153/A sky130_fd_sc_hd__a22o_1
XFILLER_38_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_46_2 dadda_fa_2_46_2/A dadda_fa_2_46_2/B dadda_fa_2_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/A dadda_fa_3_46_3/A sky130_fd_sc_hd__fa_1
XU$$4163 U$$4163/A U$$4175/B VGND VGND VPWR VPWR U$$4163/X sky130_fd_sc_hd__xor2_1
XFILLER_53_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4174 U$$4446/B1 U$$4174/A2 U$$4176/A1 U$$4174/B2 VGND VGND VPWR VPWR U$$4175/A
+ sky130_fd_sc_hd__a22o_1
XU$$3440 U$$3440/A U$$3490/B VGND VGND VPWR VPWR U$$3440/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4185 U$$4185/A U$$4197/B VGND VGND VPWR VPWR U$$4185/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_23_1 dadda_fa_5_23_1/A dadda_fa_5_23_1/B dadda_fa_5_23_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_24_0/B dadda_fa_7_23_0/A sky130_fd_sc_hd__fa_1
XU$$4196 _591_/Q U$$4196/A2 U$$4333/B1 U$$4196/B2 VGND VGND VPWR VPWR U$$4197/A sky130_fd_sc_hd__a22o_1
XU$$3451 U$$3451/A1 U$$3497/A2 U$$3453/A1 U$$3497/B2 VGND VGND VPWR VPWR U$$3452/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_39_1 U$$1548/X U$$1681/X U$$1814/X VGND VGND VPWR VPWR dadda_fa_3_40_0/CIN
+ dadda_fa_3_39_2/CIN sky130_fd_sc_hd__fa_1
XU$$3462 U$$3462/A U$$3561/A VGND VGND VPWR VPWR U$$3462/X sky130_fd_sc_hd__xor2_1
XFILLER_207_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3473 U$$4158/A1 U$$3497/A2 U$$3475/A1 U$$3497/B2 VGND VGND VPWR VPWR U$$3474/A
+ sky130_fd_sc_hd__a22o_1
XU$$3484 U$$3484/A U$$3490/B VGND VGND VPWR VPWR U$$3484/X sky130_fd_sc_hd__xor2_1
XFILLER_209_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_16_0 dadda_fa_5_16_0/A dadda_fa_5_16_0/B dadda_fa_5_16_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_17_0/A dadda_fa_6_16_0/CIN sky130_fd_sc_hd__fa_1
XU$$2750 U$$3022/B1 U$$2798/A2 U$$3024/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2751/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3495 U$$3495/A1 U$$3497/A2 U$$4045/A1 U$$3497/B2 VGND VGND VPWR VPWR U$$3496/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2761 U$$2761/A U$$2787/B VGND VGND VPWR VPWR U$$2761/X sky130_fd_sc_hd__xor2_1
XFILLER_209_1043 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2772 U$$2909/A1 U$$2814/A2 U$$2909/B1 U$$2814/B2 VGND VGND VPWR VPWR U$$2773/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2783 U$$2783/A U$$2813/B VGND VGND VPWR VPWR U$$2783/X sky130_fd_sc_hd__xor2_1
XFILLER_209_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2794 U$$4436/B1 U$$2798/A2 U$$4301/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2795/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_1118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1028 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput207 c[55] VGND VGND VPWR VPWR input207/X sky130_fd_sc_hd__clkbuf_4
XFILLER_130_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput218 c[65] VGND VGND VPWR VPWR input218/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput229 c[75] VGND VGND VPWR VPWR input229/X sky130_fd_sc_hd__clkbuf_4
XFILLER_124_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$701 final_adder.U$$701/A final_adder.U$$701/B VGND VGND VPWR VPWR
+ _247_/D sky130_fd_sc_hd__xor2_1
XFILLER_25_1042 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$712 final_adder.U$$712/A final_adder.U$$712/B VGND VGND VPWR VPWR
+ _258_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$723 final_adder.U$$723/A final_adder.U$$723/B VGND VGND VPWR VPWR
+ _269_/D sky130_fd_sc_hd__xor2_1
XTAP_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$734 ANTENNA_9/DIODE final_adder.U$$734/B VGND VGND VPWR VPWR _280_/D
+ sky130_fd_sc_hd__xor2_1
XFILLER_116_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$745 final_adder.U$$745/A final_adder.U$$745/B VGND VGND VPWR VPWR
+ _291_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_leaf_95_clk _634_/CLK VGND VGND VPWR VPWR _633_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater960 U$$3498/B VGND VGND VPWR VPWR U$$3478/B sky130_fd_sc_hd__buf_8
XU$$606 U$$880/A1 U$$616/A2 U$$745/A1 U$$616/B2 VGND VGND VPWR VPWR U$$607/A sky130_fd_sc_hd__a22o_1
Xrepeater971 U$$3423/B VGND VGND VPWR VPWR U$$3424/A sky130_fd_sc_hd__buf_8
XFILLER_44_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater982 _663_/Q VGND VGND VPWR VPWR U$$3288/A sky130_fd_sc_hd__buf_4
XU$$617 U$$617/A U$$659/B VGND VGND VPWR VPWR U$$617/X sky130_fd_sc_hd__xor2_1
XFILLER_205_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_41_1 U$$488/X U$$621/X U$$754/X VGND VGND VPWR VPWR dadda_fa_2_42_3/CIN
+ dadda_fa_2_41_5/B sky130_fd_sc_hd__fa_1
XU$$628 U$$628/A1 U$$632/A2 U$$82/A1 U$$632/B2 VGND VGND VPWR VPWR U$$629/A sky130_fd_sc_hd__a22o_1
XFILLER_72_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater993 U$$2944/B VGND VGND VPWR VPWR U$$2916/B sky130_fd_sc_hd__buf_6
XU$$639 U$$639/A U$$651/B VGND VGND VPWR VPWR U$$639/X sky130_fd_sc_hd__xor2_1
XFILLER_44_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1084 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1506 U$$4442/A1 VGND VGND VPWR VPWR U$$3346/A1 sky130_fd_sc_hd__buf_6
XFILLER_153_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1517 _575_/Q VGND VGND VPWR VPWR U$$3753/A1 sky130_fd_sc_hd__buf_6
XFILLER_126_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1528 U$$3475/B1 VGND VGND VPWR VPWR U$$600/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1539 _573_/Q VGND VGND VPWR VPWR U$$4160/A1 sky130_fd_sc_hd__buf_6
XFILLER_137_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_70_3 dadda_fa_3_70_3/A dadda_fa_3_70_3/B dadda_fa_3_70_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_1/B dadda_fa_4_70_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_63_2 dadda_fa_3_63_2/A dadda_fa_3_63_2/B dadda_fa_3_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_1/A dadda_fa_4_63_2/B sky130_fd_sc_hd__fa_1
XFILLER_0_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_56_1 dadda_fa_3_56_1/A dadda_fa_3_56_1/B dadda_fa_3_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_0/CIN dadda_fa_4_56_2/A sky130_fd_sc_hd__fa_1
XFILLER_82_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_86_clk _628_/CLK VGND VGND VPWR VPWR _626_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_33_0 dadda_fa_6_33_0/A dadda_fa_6_33_0/B dadda_fa_6_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_34_0/B dadda_fa_7_33_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_49_0 dadda_fa_3_49_0/A dadda_fa_3_49_0/B dadda_fa_3_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_0/B dadda_fa_4_49_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_207_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2002 U$$3372/A1 U$$1922/X U$$3374/A1 U$$1923/X VGND VGND VPWR VPWR U$$2003/A sky130_fd_sc_hd__a22o_1
XFILLER_74_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2013 U$$2013/A U$$2029/B VGND VGND VPWR VPWR U$$2013/X sky130_fd_sc_hd__xor2_1
XFILLER_210_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2024 U$$3255/B1 U$$2052/A2 U$$3122/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2025/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2035 U$$2035/A U$$2039/B VGND VGND VPWR VPWR U$$2035/X sky130_fd_sc_hd__xor2_1
XU$$1301 U$$614/B1 U$$1309/A2 U$$344/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1302/A sky130_fd_sc_hd__a22o_1
XU$$2046 U$$2318/B1 U$$2052/A2 U$$3418/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2047/A
+ sky130_fd_sc_hd__a22o_1
XU$$1312 U$$1312/A U$$1356/B VGND VGND VPWR VPWR U$$1312/X sky130_fd_sc_hd__xor2_1
XU$$2057 _647_/Q VGND VGND VPWR VPWR U$$2057/Y sky130_fd_sc_hd__inv_1
XU$$2068 U$$2068/A U$$2108/B VGND VGND VPWR VPWR U$$2068/X sky130_fd_sc_hd__xor2_1
XU$$1323 U$$501/A1 U$$1323/A2 U$$229/A1 U$$1323/B2 VGND VGND VPWR VPWR U$$1324/A sky130_fd_sc_hd__a22o_1
XU$$1334 U$$1334/A U$$1370/A VGND VGND VPWR VPWR U$$1334/X sky130_fd_sc_hd__xor2_1
XU$$2079 U$$981/B1 U$$2115/A2 U$$848/A1 U$$2115/B2 VGND VGND VPWR VPWR U$$2080/A sky130_fd_sc_hd__a22o_1
XFILLER_204_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1345 U$$658/B1 U$$1345/A2 U$$525/A1 U$$1345/B2 VGND VGND VPWR VPWR U$$1346/A sky130_fd_sc_hd__a22o_1
XFILLER_206_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1356 U$$1356/A U$$1356/B VGND VGND VPWR VPWR U$$1356/X sky130_fd_sc_hd__xor2_1
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_3_114_1 U$$3826/X U$$3959/X VGND VGND VPWR VPWR dadda_fa_4_115_2/B dadda_ha_3_114_1/SUM
+ sky130_fd_sc_hd__ha_1
XU$$1367 U$$817/B1 U$$1367/A2 U$$1367/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1368/A
+ sky130_fd_sc_hd__a22o_1
XU$$1378 U$$8/A1 U$$1428/A2 U$$8/B1 U$$1428/B2 VGND VGND VPWR VPWR U$$1379/A sky130_fd_sc_hd__a22o_1
XFILLER_204_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1389 U$$1389/A U$$1425/B VGND VGND VPWR VPWR U$$1389/X sky130_fd_sc_hd__xor2_1
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_106_0 dadda_fa_7_106_0/A dadda_fa_7_106_0/B dadda_fa_7_106_0/CIN VGND
+ VGND VPWR VPWR _531_/D _402_/D sky130_fd_sc_hd__fa_1
XFILLER_156_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_811 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_51_0 input203/X dadda_fa_2_51_0/B dadda_fa_2_51_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_52_0/B dadda_fa_3_51_2/B sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_77_clk _628_/CLK VGND VGND VPWR VPWR _674_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$30 _454_/Q _326_/Q VGND VGND VPWR VPWR final_adder.U$$525/B1 final_adder.U$$652/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$41 _465_/Q _337_/Q VGND VGND VPWR VPWR final_adder.U$$169/B1 final_adder.U$$663/A
+ sky130_fd_sc_hd__ha_1
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$52 _476_/Q _348_/Q VGND VGND VPWR VPWR final_adder.U$$547/B1 final_adder.U$$674/A
+ sky130_fd_sc_hd__ha_1
XFILLER_198_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3270 U$$3270/A U$$3272/B VGND VGND VPWR VPWR U$$3270/X sky130_fd_sc_hd__xor2_1
XU$$3281 U$$3281/A1 U$$3155/X U$$3283/A1 U$$3156/X VGND VGND VPWR VPWR U$$3282/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$63 _487_/Q _359_/Q VGND VGND VPWR VPWR final_adder.U$$191/B1 final_adder.U$$685/A
+ sky130_fd_sc_hd__ha_1
XU$$3292 U$$3290/Y _664_/Q _663_/Q U$$3291/X U$$3288/Y VGND VGND VPWR VPWR U$$3292/X
+ sky130_fd_sc_hd__a32o_4
Xfinal_adder.U$$74 _498_/Q _370_/Q VGND VGND VPWR VPWR final_adder.U$$569/B1 final_adder.U$$696/A
+ sky130_fd_sc_hd__ha_1
XFILLER_55_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$85 _509_/Q _381_/Q VGND VGND VPWR VPWR final_adder.U$$213/B1 final_adder.U$$707/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$96 _520_/Q _392_/Q VGND VGND VPWR VPWR final_adder.U$$591/B1 final_adder.U$$718/A
+ sky130_fd_sc_hd__ha_1
XFILLER_181_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2580 U$$2717/A1 U$$2580/A2 U$$3404/A1 U$$2580/B2 VGND VGND VPWR VPWR U$$2581/A
+ sky130_fd_sc_hd__a22o_1
XU$$2591 U$$2591/A U$$2597/B VGND VGND VPWR VPWR U$$2591/X sky130_fd_sc_hd__xor2_1
XFILLER_179_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1890 U$$1890/A U$$1917/A VGND VGND VPWR VPWR U$$1890/X sky130_fd_sc_hd__xor2_1
XFILLER_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1650_1723 VGND VGND VPWR VPWR U$$1650_1723/HI U$$1650/A1 sky130_fd_sc_hd__conb_1
XFILLER_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_80_2 dadda_fa_4_80_2/A dadda_fa_4_80_2/B dadda_fa_4_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/CIN dadda_fa_5_80_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_73_1 dadda_fa_4_73_1/A dadda_fa_4_73_1/B dadda_fa_4_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/B dadda_fa_5_73_1/B sky130_fd_sc_hd__fa_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_89_1 U$$2180/X U$$2313/X U$$2446/X VGND VGND VPWR VPWR dadda_fa_2_90_4/A
+ dadda_fa_2_89_5/B sky130_fd_sc_hd__fa_1
XFILLER_131_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_50_0 dadda_fa_7_50_0/A dadda_fa_7_50_0/B dadda_fa_7_50_0/CIN VGND VGND
+ VPWR VPWR _475_/D _346_/D sky130_fd_sc_hd__fa_2
XFILLER_135_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_66_0 dadda_fa_4_66_0/A dadda_fa_4_66_0/B dadda_fa_4_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/A dadda_fa_5_66_1/A sky130_fd_sc_hd__fa_1
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_clk _369_/CLK VGND VGND VPWR VPWR _569_/CLK sky130_fd_sc_hd__clkbuf_16
Xfinal_adder.U$$531 final_adder.U$$658/A final_adder.U$$658/B final_adder.U$$531/B1
+ VGND VGND VPWR VPWR final_adder.U$$659/B sky130_fd_sc_hd__a21o_1
XTAP_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_630_ _633_/CLK _630_/D VGND VGND VPWR VPWR _630_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$553 final_adder.U$$680/A final_adder.U$$680/B final_adder.U$$553/B1
+ VGND VGND VPWR VPWR final_adder.U$$681/B sky130_fd_sc_hd__a21o_1
XTAP_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$403 U$$403/A U$$411/A VGND VGND VPWR VPWR U$$403/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$575 final_adder.U$$702/A final_adder.U$$702/B final_adder.U$$575/B1
+ VGND VGND VPWR VPWR final_adder.U$$703/B sky130_fd_sc_hd__a21o_1
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$414 _623_/Q U$$414/B VGND VGND VPWR VPWR U$$414/X sky130_fd_sc_hd__and2_1
XFILLER_57_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$425 U$$562/A1 U$$447/A2 U$$973/B1 U$$447/B2 VGND VGND VPWR VPWR U$$426/A sky130_fd_sc_hd__a22o_1
Xrepeater790 U$$2608/X VGND VGND VPWR VPWR U$$2707/B2 sky130_fd_sc_hd__buf_6
X_561_ _569_/CLK _561_/D VGND VGND VPWR VPWR _561_/Q sky130_fd_sc_hd__dfxtp_2
Xfinal_adder.U$$597 final_adder.U$$724/A final_adder.U$$724/B final_adder.U$$597/B1
+ VGND VGND VPWR VPWR final_adder.U$$725/B sky130_fd_sc_hd__a21o_1
XFILLER_205_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$436 U$$436/A U$$532/B VGND VGND VPWR VPWR U$$436/X sky130_fd_sc_hd__xor2_1
XFILLER_84_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$447 U$$582/B1 U$$447/A2 U$$449/A1 U$$447/B2 VGND VGND VPWR VPWR U$$448/A sky130_fd_sc_hd__a22o_1
XU$$458 U$$458/A U$$536/B VGND VGND VPWR VPWR U$$458/X sky130_fd_sc_hd__xor2_1
XFILLER_189_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$469 U$$880/A1 U$$483/A2 U$$882/A1 U$$483/B2 VGND VGND VPWR VPWR U$$470/A sky130_fd_sc_hd__a22o_1
X_492_ _492_/CLK _492_/D VGND VGND VPWR VPWR _492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1303 U$$3805/B1 VGND VGND VPWR VPWR U$$4218/A1 sky130_fd_sc_hd__buf_4
Xrepeater1314 U$$3253/B1 VGND VGND VPWR VPWR U$$650/B1 sky130_fd_sc_hd__buf_4
XFILLER_153_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1325 U$$3388/B1 VGND VGND VPWR VPWR U$$785/B1 sky130_fd_sc_hd__buf_8
XFILLER_5_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1336 U$$4208/B1 VGND VGND VPWR VPWR U$$4484/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1347 U$$3519/B1 VGND VGND VPWR VPWR U$$916/B1 sky130_fd_sc_hd__buf_4
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1358 U$$4065/B1 VGND VGND VPWR VPWR U$$2832/B1 sky130_fd_sc_hd__buf_6
XFILLER_181_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1369 U$$4337/B1 VGND VGND VPWR VPWR U$$4476/A1 sky130_fd_sc_hd__buf_4
XFILLER_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_59_clk _535_/CLK VGND VGND VPWR VPWR _596_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_209_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$970 U$$970/A U$$994/B VGND VGND VPWR VPWR U$$970/X sky130_fd_sc_hd__xor2_1
XFILLER_91_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1120 U$$435/A1 U$$1150/A2 U$$985/A1 U$$1150/B2 VGND VGND VPWR VPWR U$$1121/A sky130_fd_sc_hd__a22o_1
XFILLER_62_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$981 U$$22/A1 U$$999/A2 U$$981/B1 U$$999/B2 VGND VGND VPWR VPWR U$$982/A sky130_fd_sc_hd__a22o_1
XFILLER_211_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$992 U$$992/A U$$994/B VGND VGND VPWR VPWR U$$992/X sky130_fd_sc_hd__xor2_1
XFILLER_50_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1131 U$$1131/A U$$1191/B VGND VGND VPWR VPWR U$$1131/X sky130_fd_sc_hd__xor2_1
XU$$1142 U$$2375/A1 U$$1146/A2 U$$48/A1 U$$1146/B2 VGND VGND VPWR VPWR U$$1143/A sky130_fd_sc_hd__a22o_1
XU$$1153 U$$1153/A U$$1195/B VGND VGND VPWR VPWR U$$1153/X sky130_fd_sc_hd__xor2_1
XFILLER_149_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1164 U$$68/A1 U$$1190/A2 U$$70/A1 U$$1190/B2 VGND VGND VPWR VPWR U$$1165/A sky130_fd_sc_hd__a22o_1
XFILLER_93_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1175 U$$1175/A U$$1177/B VGND VGND VPWR VPWR U$$1175/X sky130_fd_sc_hd__xor2_1
XU$$1186 U$$501/A1 U$$1208/A2 U$$229/A1 U$$1208/B2 VGND VGND VPWR VPWR U$$1187/A sky130_fd_sc_hd__a22o_1
XU$$1197 U$$1197/A U$$1203/B VGND VGND VPWR VPWR U$$1197/X sky130_fd_sc_hd__xor2_1
XFILLER_31_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_90_1 dadda_fa_5_90_1/A dadda_fa_5_90_1/B dadda_fa_5_90_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_91_0/B dadda_fa_7_90_0/A sky130_fd_sc_hd__fa_1
XFILLER_15_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_83_0 dadda_fa_5_83_0/A dadda_fa_5_83_0/B dadda_fa_5_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_84_0/A dadda_fa_6_83_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_99_0 U$$2465/Y U$$2599/X U$$2732/X VGND VGND VPWR VPWR dadda_fa_3_100_1/A
+ dadda_fa_3_99_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_75_7 U$$4413/X input229/X dadda_fa_1_75_7/CIN VGND VGND VPWR VPWR dadda_fa_2_76_2/CIN
+ dadda_fa_2_75_5/CIN sky130_fd_sc_hd__fa_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_6 dadda_fa_1_68_6/A dadda_fa_1_68_6/B dadda_fa_1_68_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_2/B dadda_fa_2_68_5/B sky130_fd_sc_hd__fa_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_109 _179_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_98_0 dadda_fa_7_98_0/A dadda_fa_7_98_0/B dadda_fa_7_98_0/CIN VGND VGND
+ VPWR VPWR _523_/D _394_/D sky130_fd_sc_hd__fa_1
XFILLER_194_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4_1760 VGND VGND VPWR VPWR U$$4_1760/HI U$$4/A3 sky130_fd_sc_hd__conb_1
Xdadda_fa_6_113_0 dadda_fa_6_113_0/A dadda_fa_6_113_0/B dadda_fa_6_113_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_114_0/B dadda_fa_7_113_0/CIN sky130_fd_sc_hd__fa_1
XTAP_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_613_ _613_/CLK _613_/D VGND VGND VPWR VPWR _613_/Q sky130_fd_sc_hd__dfxtp_2
Xfinal_adder.U$$361 final_adder.U$$360/A final_adder.U$$337/X final_adder.U$$339/X
+ VGND VGND VPWR VPWR final_adder.U$$361/X sky130_fd_sc_hd__a21o_1
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$200 U$$200/A U$$226/B VGND VGND VPWR VPWR U$$200/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$372 final_adder.U$$372/A final_adder.U$$372/B VGND VGND VPWR VPWR
+ final_adder.U$$372/X sky130_fd_sc_hd__and2_1
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$211 U$$74/A1 U$$217/A2 U$$76/A1 U$$217/B2 VGND VGND VPWR VPWR U$$212/A sky130_fd_sc_hd__a22o_1
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$383 final_adder.U$$372/X final_adder.U$$686/B final_adder.U$$373/X
+ VGND VGND VPWR VPWR final_adder.U$$718/B sky130_fd_sc_hd__a21o_2
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_33_3 dadda_fa_3_33_3/A dadda_fa_3_33_3/B dadda_fa_3_33_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_1/B dadda_fa_4_33_2/CIN sky130_fd_sc_hd__fa_1
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$222 U$$222/A U$$226/B VGND VGND VPWR VPWR U$$222/X sky130_fd_sc_hd__xor2_1
XFILLER_206_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$233 U$$96/A1 U$$249/A2 U$$98/A1 U$$249/B2 VGND VGND VPWR VPWR U$$234/A sky130_fd_sc_hd__a22o_1
XFILLER_18_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$244 U$$244/A U$$250/B VGND VGND VPWR VPWR U$$244/X sky130_fd_sc_hd__xor2_1
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_544_ _547_/CLK _544_/D VGND VGND VPWR VPWR _544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$255 U$$392/A1 U$$259/A2 U$$942/A1 U$$259/B2 VGND VGND VPWR VPWR U$$256/A sky130_fd_sc_hd__a22o_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$266 U$$266/A U$$272/B VGND VGND VPWR VPWR U$$266/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_26_2 U$$1820/B input175/X dadda_fa_3_26_2/CIN VGND VGND VPWR VPWR dadda_fa_4_27_1/A
+ dadda_fa_4_26_2/B sky130_fd_sc_hd__fa_1
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$277 _621_/Q U$$277/B VGND VGND VPWR VPWR U$$277/X sky130_fd_sc_hd__and2_1
XFILLER_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$288 U$$562/A1 U$$318/A2 U$$973/B1 U$$318/B2 VGND VGND VPWR VPWR U$$289/A sky130_fd_sc_hd__a22o_1
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$299 U$$299/A U$$309/B VGND VGND VPWR VPWR U$$299/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_19_1 U$$444/X U$$577/X U$$710/X VGND VGND VPWR VPWR dadda_fa_4_20_1/A
+ dadda_fa_4_19_2/B sky130_fd_sc_hd__fa_1
X_475_ _475_/CLK _475_/D VGND VGND VPWR VPWR _475_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1060 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$5 U$$3/B U$$5/A2 U$$1/A U$$0/Y VGND VGND VPWR VPWR U$$5/X sky130_fd_sc_hd__a22o_2
XFILLER_199_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1100 _637_/Q VGND VGND VPWR VPWR U$$1507/A sky130_fd_sc_hd__buf_4
Xrepeater1111 U$$1191/B VGND VGND VPWR VPWR U$$1151/B sky130_fd_sc_hd__buf_6
Xoutput308 _198_/Q VGND VGND VPWR VPWR o[30] sky130_fd_sc_hd__buf_2
XFILLER_142_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1122 U$$982/B VGND VGND VPWR VPWR U$$980/B sky130_fd_sc_hd__buf_6
Xoutput319 _208_/Q VGND VGND VPWR VPWR o[40] sky130_fd_sc_hd__buf_2
XFILLER_154_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1133 U$$925/B VGND VGND VPWR VPWR U$$897/B sky130_fd_sc_hd__buf_6
XFILLER_142_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1144 U$$810/B VGND VGND VPWR VPWR U$$821/A sky130_fd_sc_hd__buf_12
XU$$4471_1814 VGND VGND VPWR VPWR U$$4471_1814/HI U$$4471/B sky130_fd_sc_hd__conb_1
XFILLER_99_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1155 _625_/Q VGND VGND VPWR VPWR U$$685/A sky130_fd_sc_hd__buf_4
Xrepeater1166 U$$397/B VGND VGND VPWR VPWR U$$335/B sky130_fd_sc_hd__buf_6
XFILLER_4_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1177 U$$232/B VGND VGND VPWR VPWR U$$216/B sky130_fd_sc_hd__buf_6
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1188 U$$99/B VGND VGND VPWR VPWR U$$117/B sky130_fd_sc_hd__buf_6
Xrepeater1199 _615_/Q VGND VGND VPWR VPWR U$$956/A1 sky130_fd_sc_hd__buf_6
XFILLER_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_78_5 dadda_fa_2_78_5/A dadda_fa_2_78_5/B dadda_fa_2_78_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_2/A dadda_fa_4_78_0/A sky130_fd_sc_hd__fa_2
XFILLER_95_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3970_1758 VGND VGND VPWR VPWR U$$3970_1758/HI U$$3970/B1 sky130_fd_sc_hd__conb_1
XFILLER_208_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_970 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_811 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_108_1 dadda_fa_5_108_1/A dadda_fa_5_108_1/B dadda_fa_5_108_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_109_0/B dadda_fa_7_108_0/A sky130_fd_sc_hd__fa_2
XFILLER_144_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_80_5 U$$3093/X U$$3226/X U$$3359/X VGND VGND VPWR VPWR dadda_fa_2_81_2/B
+ dadda_fa_2_80_5/A sky130_fd_sc_hd__fa_1
XFILLER_63_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_73_4 U$$3478/X U$$3611/X U$$3744/X VGND VGND VPWR VPWR dadda_fa_2_74_1/CIN
+ dadda_fa_2_73_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_66_3 U$$3730/X U$$3863/X U$$3996/X VGND VGND VPWR VPWR dadda_fa_2_67_1/B
+ dadda_fa_2_66_4/B sky130_fd_sc_hd__fa_1
XFILLER_47_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_43_2 dadda_fa_4_43_2/A dadda_fa_4_43_2/B dadda_fa_4_43_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/CIN dadda_fa_5_43_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_59_2 U$$2386/X U$$2519/X U$$2652/X VGND VGND VPWR VPWR dadda_fa_2_60_1/A
+ dadda_fa_2_59_4/A sky130_fd_sc_hd__fa_1
XFILLER_132_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_36_1 dadda_fa_4_36_1/A dadda_fa_4_36_1/B dadda_fa_4_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/B dadda_fa_5_36_1/B sky130_fd_sc_hd__fa_1
XFILLER_6_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_13_0 dadda_fa_7_13_0/A dadda_fa_7_13_0/B dadda_fa_7_13_0/CIN VGND VGND
+ VPWR VPWR _438_/D _309_/D sky130_fd_sc_hd__fa_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1011 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_29_0 dadda_fa_4_29_0/A dadda_fa_4_29_0/B dadda_fa_4_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/A dadda_fa_5_29_1/A sky130_fd_sc_hd__fa_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_260_ _379_/CLK _260_/D VGND VGND VPWR VPWR _260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_833 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_191_ _207_/CLK _191_/D VGND VGND VPWR VPWR _191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_87 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4504 U$$4504/A1 U$$4388/X U$$4506/A1 U$$4389/X VGND VGND VPWR VPWR U$$4505/A sky130_fd_sc_hd__a22o_1
XFILLER_103_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4515 U$$4515/A U$$4515/B VGND VGND VPWR VPWR U$$4515/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_61_2 U$$927/X U$$1060/X U$$1193/X VGND VGND VPWR VPWR dadda_fa_1_62_6/B
+ dadda_fa_1_61_8/B sky130_fd_sc_hd__fa_1
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3803 U$$3803/A1 U$$3805/A2 U$$3805/A1 U$$3805/B2 VGND VGND VPWR VPWR U$$3804/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$18 U$$18/A1 U$$8/A2 U$$20/A1 U$$8/B2 VGND VGND VPWR VPWR U$$19/A sky130_fd_sc_hd__a22o_1
XU$$3814 U$$3814/A U$$3835/A VGND VGND VPWR VPWR U$$3814/X sky130_fd_sc_hd__xor2_1
XFILLER_66_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$29 U$$29/A U$$57/B VGND VGND VPWR VPWR U$$29/X sky130_fd_sc_hd__xor2_1
XFILLER_206_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3825 U$$4236/A1 U$$3833/A2 U$$4238/A1 U$$3833/B2 VGND VGND VPWR VPWR U$$3826/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3836 U$$3836/A VGND VGND VPWR VPWR U$$3836/Y sky130_fd_sc_hd__inv_1
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_0 U$$1931/X U$$2064/X input181/X VGND VGND VPWR VPWR dadda_fa_4_32_0/B
+ dadda_fa_4_31_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3847 U$$3847/A U$$3895/B VGND VGND VPWR VPWR U$$3847/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$180 final_adder.U$$675/A final_adder.U$$674/A VGND VGND VPWR VPWR
+ final_adder.U$$282/B sky130_fd_sc_hd__and2_1
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3858 U$$4269/A1 U$$3970/A2 _560_/Q U$$3970/B2 VGND VGND VPWR VPWR U$$3859/A sky130_fd_sc_hd__a22o_1
XFILLER_206_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$191 final_adder.U$$685/A final_adder.U$$557/B1 final_adder.U$$191/B1
+ VGND VGND VPWR VPWR final_adder.U$$191/X sky130_fd_sc_hd__a21o_1
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3869 U$$3869/A U$$3949/B VGND VGND VPWR VPWR U$$3869/X sky130_fd_sc_hd__xor2_1
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4429_1793 VGND VGND VPWR VPWR U$$4429_1793/HI U$$4429/B sky130_fd_sc_hd__conb_1
XFILLER_206_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_527_ _615_/CLK _527_/D VGND VGND VPWR VPWR _527_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_458_ _458_/CLK _458_/D VGND VGND VPWR VPWR _458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_389_ _520_/CLK _389_/D VGND VGND VPWR VPWR _389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_90_4 dadda_fa_2_90_4/A dadda_fa_2_90_4/B dadda_fa_2_90_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_91_1/CIN dadda_fa_3_90_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_12_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_83_3 dadda_fa_2_83_3/A dadda_fa_2_83_3/B dadda_fa_2_83_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/B dadda_fa_3_83_3/B sky130_fd_sc_hd__fa_1
XFILLER_86_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_76_2 dadda_fa_2_76_2/A dadda_fa_2_76_2/B dadda_fa_2_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/A dadda_fa_3_76_3/A sky130_fd_sc_hd__fa_1
XFILLER_141_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_53_1 dadda_fa_5_53_1/A dadda_fa_5_53_1/B dadda_fa_5_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_54_0/B dadda_fa_7_53_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_69_1 dadda_fa_2_69_1/A dadda_fa_2_69_1/B dadda_fa_2_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_0/CIN dadda_fa_3_69_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_46_0 dadda_fa_5_46_0/A dadda_fa_5_46_0/B dadda_fa_5_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_47_0/A dadda_fa_6_46_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2883_1743 VGND VGND VPWR VPWR U$$2883_1743/HI U$$2883/A1 sky130_fd_sc_hd__conb_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_831 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_120_0 U$$4503/X input152/X dadda_fa_5_120_0/CIN VGND VGND VPWR VPWR dadda_fa_6_121_0/A
+ dadda_fa_6_120_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_191_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_28 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_71_1 U$$2543/X U$$2676/X U$$2809/X VGND VGND VPWR VPWR dadda_fa_2_72_0/CIN
+ dadda_fa_2_71_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_64_0 U$$2529/X U$$2662/X U$$2795/X VGND VGND VPWR VPWR dadda_fa_2_65_0/B
+ dadda_fa_2_64_3/B sky130_fd_sc_hd__fa_1
XFILLER_87_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2409 U$$628/A1 U$$2435/A2 U$$3096/A1 U$$2435/B2 VGND VGND VPWR VPWR U$$2410/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1708 U$$3352/A1 U$$1710/A2 U$$3217/A1 U$$1710/B2 VGND VGND VPWR VPWR U$$1709/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1719 U$$1719/A U$$1719/B VGND VGND VPWR VPWR U$$1719/X sky130_fd_sc_hd__xor2_1
XFILLER_199_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_731 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_312_ _441_/CLK _312_/D VGND VGND VPWR VPWR _312_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_243_ _372_/CLK _243_/D VGND VGND VPWR VPWR _243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 a[25] VGND VGND VPWR VPWR _641_/D sky130_fd_sc_hd__clkbuf_1
X_174_ _189_/CLK _174_/D VGND VGND VPWR VPWR _174_/Q sky130_fd_sc_hd__dfxtp_1
Xinput29 a[35] VGND VGND VPWR VPWR _651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_93_2 dadda_fa_3_93_2/A dadda_fa_3_93_2/B dadda_fa_3_93_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_1/A dadda_fa_4_93_2/B sky130_fd_sc_hd__fa_1
XFILLER_202_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_86_1 dadda_fa_3_86_1/A dadda_fa_3_86_1/B dadda_fa_3_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_0/CIN dadda_fa_4_86_2/A sky130_fd_sc_hd__fa_1
XFILLER_163_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_63_0 dadda_fa_6_63_0/A dadda_fa_6_63_0/B dadda_fa_6_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_64_0/B dadda_fa_7_63_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_184_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_79_0 dadda_fa_3_79_0/A dadda_fa_3_79_0/B dadda_fa_3_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_0/B dadda_fa_4_79_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_53_0 U$$113/X U$$246/X VGND VGND VPWR VPWR dadda_fa_1_54_8/B dadda_fa_2_53_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_151_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater608 U$$219/A2 VGND VGND VPWR VPWR U$$175/A2 sky130_fd_sc_hd__buf_6
XFILLER_77_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4301 _575_/Q U$$4347/A2 U$$4301/B1 U$$4347/B2 VGND VGND VPWR VPWR U$$4302/A sky130_fd_sc_hd__a22o_1
Xrepeater619 U$$1478/A2 VGND VGND VPWR VPWR U$$1428/A2 sky130_fd_sc_hd__buf_6
XFILLER_42_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4312 U$$4312/A _679_/Q VGND VGND VPWR VPWR U$$4312/X sky130_fd_sc_hd__xor2_1
XU$$4323 U$$4323/A1 U$$4327/A2 _587_/Q U$$4333/B2 VGND VGND VPWR VPWR U$$4324/A sky130_fd_sc_hd__a22o_1
XFILLER_65_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4334 U$$4334/A U$$4334/B VGND VGND VPWR VPWR U$$4334/X sky130_fd_sc_hd__xor2_1
XU$$3600 U$$3735/B1 U$$3636/A2 U$$3602/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3601/A
+ sky130_fd_sc_hd__a22o_1
XU$$4345 U$$4482/A1 U$$4251/X U$$4484/A1 U$$4345/B2 VGND VGND VPWR VPWR U$$4346/A
+ sky130_fd_sc_hd__a22o_1
XU$$4356 U$$4356/A U$$4382/B VGND VGND VPWR VPWR U$$4356/X sky130_fd_sc_hd__xor2_1
XFILLER_93_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3611 U$$3611/A U$$3613/B VGND VGND VPWR VPWR U$$3611/X sky130_fd_sc_hd__xor2_1
XU$$3622 _578_/Q U$$3662/A2 U$$3624/A1 U$$3662/B2 VGND VGND VPWR VPWR U$$3623/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_115_1 U$$4360/X U$$4493/X input146/X VGND VGND VPWR VPWR dadda_fa_5_116_0/B
+ dadda_fa_5_115_1/B sky130_fd_sc_hd__fa_1
XU$$4367 U$$805/A1 U$$4369/A2 U$$805/B1 U$$4369/B2 VGND VGND VPWR VPWR U$$4368/A sky130_fd_sc_hd__a22o_1
XFILLER_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3633 U$$3633/A U$$3698/A VGND VGND VPWR VPWR U$$3633/X sky130_fd_sc_hd__xor2_1
XU$$4378 U$$4378/A U$$4383/A VGND VGND VPWR VPWR U$$4378/X sky130_fd_sc_hd__xor2_1
XFILLER_46_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4389 U$$4387/B U$$4384/A U$$4389/B1 U$$4384/Y VGND VGND VPWR VPWR U$$4389/X sky130_fd_sc_hd__a22o_4
XU$$3644 U$$3779/B1 U$$3674/A2 U$$3646/A1 U$$3674/B2 VGND VGND VPWR VPWR U$$3645/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3655 U$$3655/A U$$3671/B VGND VGND VPWR VPWR U$$3655/X sky130_fd_sc_hd__xor2_1
XU$$2910 U$$2910/A U$$2988/B VGND VGND VPWR VPWR U$$2910/X sky130_fd_sc_hd__xor2_1
XU$$3666 U$$3803/A1 U$$3566/X U$$3805/A1 U$$3567/X VGND VGND VPWR VPWR U$$3667/A sky130_fd_sc_hd__a22o_1
XFILLER_18_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2921 U$$3056/B1 U$$2929/A2 U$$731/A1 U$$2929/B2 VGND VGND VPWR VPWR U$$2922/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_108_0 dadda_fa_4_108_0/A dadda_fa_4_108_0/B dadda_fa_4_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/A dadda_fa_5_108_1/A sky130_fd_sc_hd__fa_1
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2932 U$$2932/A U$$2972/B VGND VGND VPWR VPWR U$$2932/X sky130_fd_sc_hd__xor2_1
XU$$3677 U$$3677/A _669_/Q VGND VGND VPWR VPWR U$$3677/X sky130_fd_sc_hd__xor2_1
XU$$3688 U$$4510/A1 U$$3688/A2 U$$4512/A1 U$$3688/B2 VGND VGND VPWR VPWR U$$3689/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_399 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2943 U$$3626/B1 U$$2943/A2 U$$3493/A1 U$$2943/B2 VGND VGND VPWR VPWR U$$2944/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2954 U$$2954/A U$$2988/B VGND VGND VPWR VPWR U$$2954/X sky130_fd_sc_hd__xor2_1
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3699 U$$3699/A VGND VGND VPWR VPWR U$$3699/Y sky130_fd_sc_hd__inv_1
XU$$2965 U$$4333/B1 U$$2981/A2 U$$4198/B1 U$$2981/B2 VGND VGND VPWR VPWR U$$2966/A
+ sky130_fd_sc_hd__a22o_1
XU$$2976 U$$2976/A U$$3008/B VGND VGND VPWR VPWR U$$2976/X sky130_fd_sc_hd__xor2_1
XU$$2987 U$$3124/A1 U$$2997/A2 U$$3124/B1 U$$2997/B2 VGND VGND VPWR VPWR U$$2988/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_270 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_281 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2998 U$$2998/A U$$3000/B VGND VGND VPWR VPWR U$$2998/X sky130_fd_sc_hd__xor2_1
XFILLER_34_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_438 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_292 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_81_0 U$$4425/X input236/X dadda_fa_2_81_0/CIN VGND VGND VPWR VPWR dadda_fa_3_82_0/B
+ dadda_fa_3_81_2/B sky130_fd_sc_hd__fa_1
Xdadda_ha_1_51_8 U$$3301/X U$$3434/X VGND VGND VPWR VPWR dadda_fa_2_52_3/A dadda_fa_3_51_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_103_917 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_50_6 U$$2501/X U$$2634/X U$$2767/X VGND VGND VPWR VPWR dadda_fa_2_51_2/B
+ dadda_fa_2_50_5/B sky130_fd_sc_hd__fa_1
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_2_0 U$$180/B input179/X dadda_ha_6_2_0/SUM VGND VGND VPWR VPWR _427_/D
+ _298_/D sky130_fd_sc_hd__fa_1
XFILLER_52_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1039 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_950 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_80_0 dadda_fa_7_80_0/A dadda_fa_7_80_0/B dadda_fa_7_80_0/CIN VGND VGND
+ VPWR VPWR _505_/D _376_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_96_0 dadda_fa_4_96_0/A dadda_fa_4_96_0/B dadda_fa_4_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/A dadda_fa_5_96_1/A sky130_fd_sc_hd__fa_1
XFILLER_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2206 U$$2343/A1 U$$2242/A2 U$$2345/A1 U$$2242/B2 VGND VGND VPWR VPWR U$$2207/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2217 U$$2217/A U$$2263/B VGND VGND VPWR VPWR U$$2217/X sky130_fd_sc_hd__xor2_1
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2228 U$$310/A1 U$$2248/A2 U$$584/B1 U$$2248/B2 VGND VGND VPWR VPWR U$$2229/A sky130_fd_sc_hd__a22o_1
XU$$2239 U$$2239/A U$$2241/B VGND VGND VPWR VPWR U$$2239/X sky130_fd_sc_hd__xor2_1
XFILLER_16_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1505 U$$1505/A U$$1507/A VGND VGND VPWR VPWR U$$1505/X sky130_fd_sc_hd__xor2_1
XFILLER_63_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1516 U$$1516/A U$$1558/B VGND VGND VPWR VPWR U$$1516/X sky130_fd_sc_hd__xor2_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1527 U$$705/A1 U$$1553/A2 U$$568/B1 U$$1553/B2 VGND VGND VPWR VPWR U$$1528/A sky130_fd_sc_hd__a22o_1
XU$$1538 U$$1538/A U$$1578/B VGND VGND VPWR VPWR U$$1538/X sky130_fd_sc_hd__xor2_1
XFILLER_167_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1549 U$$999/B1 U$$1561/A2 U$$866/A1 U$$1561/B2 VGND VGND VPWR VPWR U$$1550/A sky130_fd_sc_hd__a22o_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_226_ _353_/CLK _226_/D VGND VGND VPWR VPWR _226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_959 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_5 dadda_fa_2_60_5/A dadda_fa_2_60_5/B dadda_fa_2_60_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_2/A dadda_fa_4_60_0/A sky130_fd_sc_hd__fa_2
Xrepeater405 U$$795/A2 VGND VGND VPWR VPWR U$$725/A2 sky130_fd_sc_hd__buf_4
Xrepeater416 U$$552/X VGND VGND VPWR VPWR U$$668/A2 sky130_fd_sc_hd__buf_4
Xrepeater427 U$$491/A2 VGND VGND VPWR VPWR U$$499/A2 sky130_fd_sc_hd__buf_6
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_53_4 dadda_fa_2_53_4/A dadda_fa_2_53_4/B dadda_fa_2_53_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/CIN dadda_fa_3_53_3/CIN sky130_fd_sc_hd__fa_1
XU$$4120 U$$4394/A1 U$$4140/A2 U$$4396/A1 U$$4140/B2 VGND VGND VPWR VPWR U$$4121/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater438 U$$4114/X VGND VGND VPWR VPWR U$$4202/A2 sky130_fd_sc_hd__buf_6
Xrepeater449 U$$4071/A2 VGND VGND VPWR VPWR U$$4061/A2 sky130_fd_sc_hd__buf_4
XFILLER_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4131 U$$4131/A U$$4215/B VGND VGND VPWR VPWR U$$4131/X sky130_fd_sc_hd__xor2_1
XU$$4142 U$$4416/A1 U$$4182/A2 U$$4418/A1 U$$4182/B2 VGND VGND VPWR VPWR U$$4143/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4153 U$$4153/A U$$4183/B VGND VGND VPWR VPWR U$$4153/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_46_3 dadda_fa_2_46_3/A dadda_fa_2_46_3/B dadda_fa_2_46_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/B dadda_fa_3_46_3/B sky130_fd_sc_hd__fa_1
XFILLER_38_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4164 _575_/Q U$$4174/A2 U$$4440/A1 U$$4174/B2 VGND VGND VPWR VPWR U$$4165/A sky130_fd_sc_hd__a22o_1
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3430 U$$3428/B U$$3425/A _666_/Q U$$3425/Y VGND VGND VPWR VPWR U$$3430/X sky130_fd_sc_hd__a22o_4
XU$$4175 U$$4175/A U$$4175/B VGND VGND VPWR VPWR U$$4175/X sky130_fd_sc_hd__xor2_1
XU$$4186 U$$4186/A1 U$$4196/A2 _587_/Q U$$4196/B2 VGND VGND VPWR VPWR U$$4187/A sky130_fd_sc_hd__a22o_1
XU$$3441 U$$3578/A1 U$$3519/A2 U$$3578/B1 U$$3519/B2 VGND VGND VPWR VPWR U$$3442/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4197 U$$4197/A U$$4197/B VGND VGND VPWR VPWR U$$4197/X sky130_fd_sc_hd__xor2_1
XU$$3452 U$$3452/A U$$3498/B VGND VGND VPWR VPWR U$$3452/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3463 U$$3735/B1 U$$3559/A2 U$$3602/A1 U$$3559/B2 VGND VGND VPWR VPWR U$$3464/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_39_2 U$$1947/X U$$2080/X U$$2213/X VGND VGND VPWR VPWR dadda_fa_3_40_1/A
+ dadda_fa_3_39_3/A sky130_fd_sc_hd__fa_1
XU$$3474 U$$3474/A U$$3498/B VGND VGND VPWR VPWR U$$3474/X sky130_fd_sc_hd__xor2_1
XFILLER_207_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3485 U$$3485/A1 U$$3519/A2 U$$3624/A1 U$$3519/B2 VGND VGND VPWR VPWR U$$3486/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_16_1 dadda_fa_5_16_1/A dadda_fa_5_16_1/B dadda_fa_5_16_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_17_0/B dadda_fa_7_16_0/A sky130_fd_sc_hd__fa_1
XU$$2740 _655_/Q VGND VGND VPWR VPWR U$$2740/Y sky130_fd_sc_hd__inv_1
XU$$2751 U$$2751/A U$$2795/B VGND VGND VPWR VPWR U$$2751/X sky130_fd_sc_hd__xor2_1
XU$$3496 U$$3496/A U$$3498/B VGND VGND VPWR VPWR U$$3496/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2762 U$$3310/A1 U$$2812/A2 U$$3447/B1 U$$2812/B2 VGND VGND VPWR VPWR U$$2763/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2773 U$$2773/A U$$2827/B VGND VGND VPWR VPWR U$$2773/X sky130_fd_sc_hd__xor2_1
XFILLER_209_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2784 U$$3056/B1 U$$2788/A2 U$$866/B1 U$$2788/B2 VGND VGND VPWR VPWR U$$2785/A
+ sky130_fd_sc_hd__a22o_1
XU$$2795 U$$2795/A U$$2795/B VGND VGND VPWR VPWR U$$2795/X sky130_fd_sc_hd__xor2_1
XFILLER_33_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1015 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_861 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_1_42_4 U$$1687/X U$$1820/X VGND VGND VPWR VPWR dadda_fa_2_43_4/B dadda_fa_3_42_0/A
+ sky130_fd_sc_hd__ha_1
Xinput208 c[56] VGND VGND VPWR VPWR input208/X sky130_fd_sc_hd__clkbuf_4
Xinput219 c[66] VGND VGND VPWR VPWR input219/X sky130_fd_sc_hd__clkbuf_1
XTAP_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$702 final_adder.U$$702/A final_adder.U$$702/B VGND VGND VPWR VPWR
+ _248_/D sky130_fd_sc_hd__xor2_1
XTAP_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$713 final_adder.U$$713/A final_adder.U$$713/B VGND VGND VPWR VPWR
+ _259_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$724 final_adder.U$$724/A final_adder.U$$724/B VGND VGND VPWR VPWR
+ _270_/D sky130_fd_sc_hd__xor2_1
XFILLER_25_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_4_12_2 U$$829/X U$$859/B VGND VGND VPWR VPWR dadda_fa_5_13_0/CIN dadda_ha_4_12_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_84_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$735 final_adder.U$$735/A final_adder.U$$735/B VGND VGND VPWR VPWR
+ _281_/D sky130_fd_sc_hd__xor2_4
Xfinal_adder.U$$746 final_adder.U$$746/A final_adder.U$$746/B VGND VGND VPWR VPWR
+ _292_/D sky130_fd_sc_hd__xor2_4
Xrepeater950 U$$3698/A VGND VGND VPWR VPWR U$$3637/B sky130_fd_sc_hd__buf_12
Xrepeater961 U$$3562/A VGND VGND VPWR VPWR U$$3498/B sky130_fd_sc_hd__buf_8
XU$$607 U$$607/A U$$613/B VGND VGND VPWR VPWR U$$607/X sky130_fd_sc_hd__xor2_1
XFILLER_29_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater972 U$$3425/A VGND VGND VPWR VPWR U$$3423/B sky130_fd_sc_hd__buf_4
XFILLER_186_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$618 U$$890/B1 U$$632/A2 U$$757/A1 U$$632/B2 VGND VGND VPWR VPWR U$$619/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_41_2 U$$887/X U$$1020/X U$$1153/X VGND VGND VPWR VPWR dadda_fa_2_42_4/A
+ dadda_fa_2_41_5/CIN sky130_fd_sc_hd__fa_2
Xrepeater983 _663_/Q VGND VGND VPWR VPWR U$$3276/B sky130_fd_sc_hd__buf_6
XFILLER_99_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$629 U$$629/A U$$659/B VGND VGND VPWR VPWR U$$629/X sky130_fd_sc_hd__xor2_1
Xrepeater994 U$$2966/B VGND VGND VPWR VPWR U$$2944/B sky130_fd_sc_hd__buf_8
XFILLER_147_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_11_0 U$$29/X U$$162/X U$$295/X VGND VGND VPWR VPWR dadda_fa_5_12_0/B dadda_fa_5_11_1/B
+ sky130_fd_sc_hd__fa_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_892 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1507 _577_/Q VGND VGND VPWR VPWR U$$4442/A1 sky130_fd_sc_hd__buf_6
XFILLER_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_115_0 U$$3561/Y U$$3695/X U$$3828/X VGND VGND VPWR VPWR dadda_fa_4_116_2/B
+ dadda_fa_4_115_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater1518 U$$52/B1 VGND VGND VPWR VPWR U$$876/A1 sky130_fd_sc_hd__buf_4
XFILLER_152_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1529 U$$3475/B1 VGND VGND VPWR VPWR U$$52/A1 sky130_fd_sc_hd__buf_8
XFILLER_153_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_63_3 dadda_fa_3_63_3/A dadda_fa_3_63_3/B dadda_fa_3_63_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_1/B dadda_fa_4_63_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_56_2 dadda_fa_3_56_2/A dadda_fa_3_56_2/B dadda_fa_3_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_1/A dadda_fa_4_56_2/B sky130_fd_sc_hd__fa_1
XFILLER_0_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_49_1 dadda_fa_3_49_1/A dadda_fa_3_49_1/B dadda_fa_3_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_0/CIN dadda_fa_4_49_2/A sky130_fd_sc_hd__fa_1
XFILLER_207_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_26_0 dadda_fa_6_26_0/A dadda_fa_6_26_0/B dadda_fa_6_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_27_0/B dadda_fa_7_26_0/CIN sky130_fd_sc_hd__fa_1
XU$$2003 U$$2003/A U$$2003/B VGND VGND VPWR VPWR U$$2003/X sky130_fd_sc_hd__xor2_1
XFILLER_62_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_528 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2014 U$$916/B1 U$$2028/A2 U$$98/A1 U$$2028/B2 VGND VGND VPWR VPWR U$$2015/A sky130_fd_sc_hd__a22o_1
XU$$2025 U$$2025/A U$$2054/A VGND VGND VPWR VPWR U$$2025/X sky130_fd_sc_hd__xor2_1
XFILLER_210_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2036 U$$940/A1 U$$2038/A2 U$$940/B1 U$$2038/B2 VGND VGND VPWR VPWR U$$2037/A sky130_fd_sc_hd__a22o_1
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1302 U$$1302/A U$$1310/B VGND VGND VPWR VPWR U$$1302/X sky130_fd_sc_hd__xor2_1
XU$$2047 U$$2047/A U$$2054/A VGND VGND VPWR VPWR U$$2047/X sky130_fd_sc_hd__xor2_1
XU$$1313 U$$2957/A1 U$$1355/A2 U$$80/B1 U$$1355/B2 VGND VGND VPWR VPWR U$$1314/A sky130_fd_sc_hd__a22o_1
XFILLER_188_500 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2058 U$$2174/B U$$2058/B VGND VGND VPWR VPWR U$$2058/X sky130_fd_sc_hd__and2_1
XU$$2069 U$$2343/A1 U$$2109/A2 U$$2345/A1 U$$2109/B2 VGND VGND VPWR VPWR U$$2070/A
+ sky130_fd_sc_hd__a22o_1
XU$$1324 U$$1324/A U$$1332/B VGND VGND VPWR VPWR U$$1324/X sky130_fd_sc_hd__xor2_1
XFILLER_167_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1335 U$$2705/A1 U$$1237/X U$$926/A1 U$$1238/X VGND VGND VPWR VPWR U$$1336/A sky130_fd_sc_hd__a22o_1
XFILLER_43_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1346 U$$1346/A U$$1369/A VGND VGND VPWR VPWR U$$1346/X sky130_fd_sc_hd__xor2_1
XFILLER_206_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1357 U$$2588/B1 U$$1367/A2 U$$948/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1358/A
+ sky130_fd_sc_hd__a22o_1
XU$$1368 U$$1368/A U$$1368/B VGND VGND VPWR VPWR U$$1368/X sky130_fd_sc_hd__xor2_1
XFILLER_204_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1379 U$$1379/A U$$1429/B VGND VGND VPWR VPWR U$$1379/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_209_ _213_/CLK _209_/D VGND VGND VPWR VPWR _209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_861 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_51_1 dadda_fa_2_51_1/A dadda_fa_2_51_1/B dadda_fa_2_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_0/CIN dadda_fa_3_51_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_44_0 U$$2356/X U$$2489/X U$$2622/X VGND VGND VPWR VPWR dadda_fa_3_45_0/B
+ dadda_fa_3_44_2/B sky130_fd_sc_hd__fa_1
XFILLER_26_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$20 _444_/Q _316_/Q VGND VGND VPWR VPWR final_adder.U$$515/B1 final_adder.U$$642/A
+ sky130_fd_sc_hd__ha_2
XU$$3260 U$$3260/A U$$3272/B VGND VGND VPWR VPWR U$$3260/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$31 _455_/Q _327_/Q VGND VGND VPWR VPWR final_adder.U$$159/B1 final_adder.U$$653/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$42 _466_/Q _338_/Q VGND VGND VPWR VPWR final_adder.U$$537/B1 final_adder.U$$664/A
+ sky130_fd_sc_hd__ha_1
XU$$3271 U$$940/B1 U$$3273/A2 U$$3273/A1 U$$3273/B2 VGND VGND VPWR VPWR U$$3272/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$53 _477_/Q _349_/Q VGND VGND VPWR VPWR final_adder.U$$181/B1 final_adder.U$$675/A
+ sky130_fd_sc_hd__ha_1
XFILLER_59_1150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3282 U$$3282/A U$$3288/A VGND VGND VPWR VPWR U$$3282/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$64 _488_/Q _360_/Q VGND VGND VPWR VPWR final_adder.U$$559/B1 final_adder.U$$686/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$75 _499_/Q _371_/Q VGND VGND VPWR VPWR final_adder.U$$203/B1 final_adder.U$$697/A
+ sky130_fd_sc_hd__ha_1
XU$$3293 U$$3291/B _663_/Q _664_/Q U$$3288/Y VGND VGND VPWR VPWR U$$3293/X sky130_fd_sc_hd__a22o_4
Xfinal_adder.U$$86 _510_/Q _382_/Q VGND VGND VPWR VPWR final_adder.U$$581/B1 final_adder.U$$708/A
+ sky130_fd_sc_hd__ha_1
XU$$2570 U$$4214/A1 U$$2470/X U$$4353/A1 U$$2471/X VGND VGND VPWR VPWR U$$2571/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$97 _521_/Q _393_/Q VGND VGND VPWR VPWR final_adder.U$$225/B1 final_adder.U$$719/A
+ sky130_fd_sc_hd__ha_1
XFILLER_185_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2581 U$$2581/A U$$2583/B VGND VGND VPWR VPWR U$$2581/X sky130_fd_sc_hd__xor2_1
XU$$2592 _611_/Q U$$2600/A2 _612_/Q U$$2600/B2 VGND VGND VPWR VPWR U$$2593/A sky130_fd_sc_hd__a22o_1
XFILLER_181_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1880 U$$1880/A U$$1884/B VGND VGND VPWR VPWR U$$1880/X sky130_fd_sc_hd__xor2_1
XFILLER_194_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1891 U$$3124/A1 U$$1897/A2 U$$3124/B1 U$$1897/B2 VGND VGND VPWR VPWR U$$1892/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_73_2 dadda_fa_4_73_2/A dadda_fa_4_73_2/B dadda_fa_4_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/CIN dadda_fa_5_73_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_157_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_89_2 U$$2579/X U$$2712/X U$$2845/X VGND VGND VPWR VPWR dadda_fa_2_90_4/B
+ dadda_fa_2_89_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_66_1 dadda_fa_4_66_1/A dadda_fa_4_66_1/B dadda_fa_4_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/B dadda_fa_5_66_1/B sky130_fd_sc_hd__fa_1
XTAP_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_43_0 dadda_fa_7_43_0/A dadda_fa_7_43_0/B dadda_fa_7_43_0/CIN VGND VGND
+ VPWR VPWR _468_/D _339_/D sky130_fd_sc_hd__fa_2
XTAP_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_59_0 dadda_fa_4_59_0/A dadda_fa_4_59_0/B dadda_fa_4_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/A dadda_fa_5_59_1/A sky130_fd_sc_hd__fa_1
XFILLER_131_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$521 final_adder.U$$648/A final_adder.U$$648/B final_adder.U$$521/B1
+ VGND VGND VPWR VPWR final_adder.U$$649/B sky130_fd_sc_hd__a21o_1
XTAP_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$543 final_adder.U$$670/A final_adder.U$$670/B final_adder.U$$543/B1
+ VGND VGND VPWR VPWR final_adder.U$$671/B sky130_fd_sc_hd__a21o_1
XFILLER_151_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_55 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$404 U$$676/B1 U$$408/A2 U$$406/A1 U$$408/B2 VGND VGND VPWR VPWR U$$405/A sky130_fd_sc_hd__a22o_1
XFILLER_56_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$565 final_adder.U$$692/A final_adder.U$$692/B final_adder.U$$565/B1
+ VGND VGND VPWR VPWR final_adder.U$$693/B sky130_fd_sc_hd__a21o_1
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater780 U$$2866/B2 VGND VGND VPWR VPWR U$$2856/B2 sky130_fd_sc_hd__buf_4
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$415 U$$413/Y _622_/Q U$$411/A U$$414/X U$$411/Y VGND VGND VPWR VPWR U$$415/X sky130_fd_sc_hd__a32o_4
XFILLER_72_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_560_ _560_/CLK _560_/D VGND VGND VPWR VPWR _560_/Q sky130_fd_sc_hd__dfxtp_4
Xfinal_adder.U$$587 final_adder.U$$714/A final_adder.U$$714/B final_adder.U$$587/B1
+ VGND VGND VPWR VPWR final_adder.U$$715/B sky130_fd_sc_hd__a21o_1
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater791 U$$2566/B2 VGND VGND VPWR VPWR U$$2550/B2 sky130_fd_sc_hd__buf_4
XFILLER_57_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$426 U$$426/A U$$456/B VGND VGND VPWR VPWR U$$426/X sky130_fd_sc_hd__xor2_1
XFILLER_72_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$437 U$$26/A1 U$$457/A2 U$$28/A1 U$$457/B2 VGND VGND VPWR VPWR U$$438/A sky130_fd_sc_hd__a22o_1
XFILLER_45_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$448 U$$448/A U$$452/B VGND VGND VPWR VPWR U$$448/X sky130_fd_sc_hd__xor2_1
XU$$459 U$$596/A1 U$$491/A2 U$$596/B1 U$$491/B2 VGND VGND VPWR VPWR U$$460/A sky130_fd_sc_hd__a22o_1
X_491_ _491_/CLK _491_/D VGND VGND VPWR VPWR _491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1304 U$$3805/B1 VGND VGND VPWR VPWR U$$2983/B1 sky130_fd_sc_hd__buf_8
Xrepeater1315 U$$2431/B1 VGND VGND VPWR VPWR U$$924/B1 sky130_fd_sc_hd__buf_6
Xrepeater1326 _599_/Q VGND VGND VPWR VPWR U$$3388/B1 sky130_fd_sc_hd__buf_4
XFILLER_165_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1337 U$$3934/B1 VGND VGND VPWR VPWR U$$4208/B1 sky130_fd_sc_hd__buf_6
Xrepeater1348 U$$3658/A1 VGND VGND VPWR VPWR U$$3519/B1 sky130_fd_sc_hd__buf_4
XFILLER_5_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1359 U$$4065/B1 VGND VGND VPWR VPWR U$$368/A1 sky130_fd_sc_hd__buf_6
XFILLER_113_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_498 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_61_0 dadda_fa_3_61_0/A dadda_fa_3_61_0/B dadda_fa_3_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_0/B dadda_fa_4_61_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_77_0 U$$958/Y U$$1092/X U$$1225/X VGND VGND VPWR VPWR dadda_fa_1_78_8/CIN
+ dadda_fa_2_77_0/A sky130_fd_sc_hd__fa_2
XFILLER_94_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$960 _630_/Q VGND VGND VPWR VPWR U$$962/B sky130_fd_sc_hd__inv_1
Xdadda_ha_4_8_0 U$$23/X U$$156/X VGND VGND VPWR VPWR dadda_fa_5_9_1/B dadda_ha_4_8_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$1110 U$$14/A1 U$$1146/A2 U$$16/A1 U$$1146/B2 VGND VGND VPWR VPWR U$$1111/A sky130_fd_sc_hd__a22o_1
XU$$971 U$$971/A1 U$$995/A2 U$$973/A1 U$$995/B2 VGND VGND VPWR VPWR U$$972/A sky130_fd_sc_hd__a22o_1
XU$$1121 U$$1121/A U$$1151/B VGND VGND VPWR VPWR U$$1121/X sky130_fd_sc_hd__xor2_1
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$982 U$$982/A U$$982/B VGND VGND VPWR VPWR U$$982/X sky130_fd_sc_hd__xor2_1
XFILLER_204_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1132 U$$719/B1 U$$1150/A2 U$$997/A1 U$$1150/B2 VGND VGND VPWR VPWR U$$1133/A sky130_fd_sc_hd__a22o_1
XFILLER_189_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$993 U$$993/A1 U$$995/A2 U$$36/A1 U$$995/B2 VGND VGND VPWR VPWR U$$994/A sky130_fd_sc_hd__a22o_1
XU$$1143 U$$1143/A U$$1147/B VGND VGND VPWR VPWR U$$1143/X sky130_fd_sc_hd__xor2_1
XFILLER_16_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1154 U$$58/A1 U$$1194/A2 U$$60/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1155/A sky130_fd_sc_hd__a22o_1
XFILLER_50_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1165 U$$1165/A U$$1191/B VGND VGND VPWR VPWR U$$1165/X sky130_fd_sc_hd__xor2_1
XFILLER_203_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1176 U$$80/A1 U$$1176/A2 U$$80/B1 U$$1176/B2 VGND VGND VPWR VPWR U$$1177/A sky130_fd_sc_hd__a22o_1
XFILLER_189_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1187 U$$1187/A U$$1209/B VGND VGND VPWR VPWR U$$1187/X sky130_fd_sc_hd__xor2_1
XU$$1198 U$$2705/A1 U$$1208/A2 U$$926/A1 U$$1208/B2 VGND VGND VPWR VPWR U$$1199/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_782 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_731 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1056 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_83_1 dadda_fa_5_83_1/A dadda_fa_5_83_1/B dadda_fa_5_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_84_0/B dadda_fa_7_83_0/A sky130_fd_sc_hd__fa_2
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_99_1 U$$2865/X U$$2998/X U$$3131/X VGND VGND VPWR VPWR dadda_fa_3_100_1/B
+ dadda_fa_3_99_3/A sky130_fd_sc_hd__fa_1
XFILLER_132_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_76_0 dadda_fa_5_76_0/A dadda_fa_5_76_0/B dadda_fa_5_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_77_0/A dadda_fa_6_76_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_75_8 dadda_fa_1_75_8/A dadda_fa_1_75_8/B dadda_fa_1_75_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_76_3/A dadda_fa_3_75_0/A sky130_fd_sc_hd__fa_2
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_7 dadda_fa_1_68_7/A dadda_fa_1_68_7/B dadda_fa_1_68_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_2/CIN dadda_fa_2_68_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_85_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_973 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3090 U$$3362/B1 U$$3110/A2 U$$4051/A1 U$$3110/B2 VGND VGND VPWR VPWR U$$3091/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_94_0 dadda_fa_1_94_0/A U$$2190/X U$$2323/X VGND VGND VPWR VPWR dadda_fa_2_95_5/B
+ dadda_fa_2_94_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_200_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$340 final_adder.U$$340/A final_adder.U$$340/B VGND VGND VPWR VPWR
+ final_adder.U$$362/B sky130_fd_sc_hd__and2_1
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$362 final_adder.U$$362/A final_adder.U$$362/B VGND VGND VPWR VPWR
+ final_adder.U$$372/A sky130_fd_sc_hd__and2_1
X_612_ _613_/CLK _612_/D VGND VGND VPWR VPWR _612_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$201 U$$201/A1 U$$219/A2 U$$749/B1 U$$219/B2 VGND VGND VPWR VPWR U$$202/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_106_0 dadda_fa_6_106_0/A dadda_fa_6_106_0/B dadda_fa_6_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_107_0/B dadda_fa_7_106_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$373 final_adder.U$$372/A final_adder.U$$361/X final_adder.U$$363/X
+ VGND VGND VPWR VPWR final_adder.U$$373/X sky130_fd_sc_hd__a21o_1
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$212 U$$212/A U$$216/B VGND VGND VPWR VPWR U$$212/X sky130_fd_sc_hd__xor2_1
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$223 U$$86/A1 U$$263/A2 U$$88/A1 U$$263/B2 VGND VGND VPWR VPWR U$$224/A sky130_fd_sc_hd__a22o_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$395 final_adder.U$$358/B final_adder.U$$670/B final_adder.U$$333/X
+ VGND VGND VPWR VPWR final_adder.U$$678/B sky130_fd_sc_hd__a21o_1
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$234 U$$234/A U$$250/B VGND VGND VPWR VPWR U$$234/X sky130_fd_sc_hd__xor2_1
XFILLER_206_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$245 U$$517/B1 U$$249/A2 U$$382/B1 U$$249/B2 VGND VGND VPWR VPWR U$$246/A sky130_fd_sc_hd__a22o_1
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_543_ _547_/CLK _543_/D VGND VGND VPWR VPWR _543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$256 U$$256/A U$$264/B VGND VGND VPWR VPWR U$$256/X sky130_fd_sc_hd__xor2_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_26_3 dadda_fa_3_26_3/A dadda_fa_3_26_3/B dadda_fa_3_26_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_27_1/B dadda_fa_4_26_2/CIN sky130_fd_sc_hd__fa_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$267 U$$676/B1 U$$141/X U$$406/A1 U$$142/X VGND VGND VPWR VPWR U$$268/A sky130_fd_sc_hd__a22o_1
XU$$278 U$$276/Y _620_/Q _619_/Q U$$277/X U$$274/Y VGND VGND VPWR VPWR U$$278/X sky130_fd_sc_hd__a32o_1
XFILLER_55_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$289 U$$289/A U$$309/B VGND VGND VPWR VPWR U$$289/X sky130_fd_sc_hd__xor2_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_474_ _475_/CLK _474_/D VGND VGND VPWR VPWR _474_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_93_0 dadda_fa_6_93_0/A dadda_fa_6_93_0/B dadda_fa_6_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_94_0/B dadda_fa_7_93_0/CIN sky130_fd_sc_hd__fa_1
XU$$6 U$$6/A1 U$$8/A2 U$$8/A1 U$$8/B2 VGND VGND VPWR VPWR U$$7/A sky130_fd_sc_hd__a22o_1
Xrepeater1101 U$$1369/A VGND VGND VPWR VPWR U$$1356/B sky130_fd_sc_hd__buf_8
XFILLER_138_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1112 U$$1177/B VGND VGND VPWR VPWR U$$1147/B sky130_fd_sc_hd__buf_6
XFILLER_5_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_444 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput309 _199_/Q VGND VGND VPWR VPWR o[31] sky130_fd_sc_hd__buf_2
XFILLER_153_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1123 U$$982/B VGND VGND VPWR VPWR U$$1040/B sky130_fd_sc_hd__buf_6
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1134 U$$951/B VGND VGND VPWR VPWR U$$925/B sky130_fd_sc_hd__buf_8
Xrepeater1145 U$$804/B VGND VGND VPWR VPWR U$$810/B sky130_fd_sc_hd__buf_12
XFILLER_154_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1156 U$$536/B VGND VGND VPWR VPWR U$$456/B sky130_fd_sc_hd__buf_6
XFILLER_99_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1167 U$$411/A VGND VGND VPWR VPWR U$$397/B sky130_fd_sc_hd__buf_6
XFILLER_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1178 U$$232/B VGND VGND VPWR VPWR U$$250/B sky130_fd_sc_hd__buf_6
XFILLER_206_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1189 U$$129/B VGND VGND VPWR VPWR U$$99/B sky130_fd_sc_hd__buf_12
XFILLER_136_1130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1090 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$790 U$$790/A U$$810/B VGND VGND VPWR VPWR U$$790/X sky130_fd_sc_hd__xor2_1
XFILLER_35_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_982 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_80_6 U$$3492/X U$$3625/X U$$3758/X VGND VGND VPWR VPWR dadda_fa_2_81_2/CIN
+ dadda_fa_2_80_5/B sky130_fd_sc_hd__fa_1
Xrepeater1690 U$$3024/B1 VGND VGND VPWR VPWR U$$2613/B1 sky130_fd_sc_hd__buf_6
XFILLER_113_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_73_5 U$$3877/X U$$4010/X U$$4143/X VGND VGND VPWR VPWR dadda_fa_2_74_2/A
+ dadda_fa_2_73_5/A sky130_fd_sc_hd__fa_1
XFILLER_141_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4487_1822 VGND VGND VPWR VPWR U$$4487_1822/HI U$$4487/B sky130_fd_sc_hd__conb_1
Xdadda_fa_1_66_4 U$$4129/X U$$4262/X U$$4395/X VGND VGND VPWR VPWR dadda_fa_2_67_1/CIN
+ dadda_fa_2_66_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_59_3 U$$2785/X U$$2918/X U$$3051/X VGND VGND VPWR VPWR dadda_fa_2_60_1/B
+ dadda_fa_2_59_4/B sky130_fd_sc_hd__fa_1
XFILLER_132_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_36_2 dadda_fa_4_36_2/A dadda_fa_4_36_2/B dadda_fa_4_36_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/CIN dadda_fa_5_36_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_1023 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_29_1 dadda_fa_4_29_1/A dadda_fa_4_29_1/B dadda_fa_4_29_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/B dadda_fa_5_29_1/B sky130_fd_sc_hd__fa_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_190_ _207_/CLK _190_/D VGND VGND VPWR VPWR _190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_62_5 U$$2126/X U$$2259/X VGND VGND VPWR VPWR dadda_fa_1_63_7/A dadda_fa_2_62_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4505 U$$4505/A U$$4505/B VGND VGND VPWR VPWR U$$4505/X sky130_fd_sc_hd__xor2_1
XU$$4516 U$$4516/A1 U$$4388/X U$$4516/B1 U$$4516/B2 VGND VGND VPWR VPWR U$$4517/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_61_3 U$$1326/X U$$1459/X U$$1592/X VGND VGND VPWR VPWR dadda_fa_1_62_6/CIN
+ dadda_fa_1_61_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$19 U$$19/A U$$9/B VGND VGND VPWR VPWR U$$19/X sky130_fd_sc_hd__xor2_1
XFILLER_18_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3804 U$$3804/A U$$3804/B VGND VGND VPWR VPWR U$$3804/X sky130_fd_sc_hd__xor2_1
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3815 U$$4361/B1 U$$3823/A2 U$$4502/A1 U$$3823/B2 VGND VGND VPWR VPWR U$$3816/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3826 U$$3826/A U$$3832/B VGND VGND VPWR VPWR U$$3826/X sky130_fd_sc_hd__xor2_1
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3837 _672_/Q VGND VGND VPWR VPWR U$$3839/B sky130_fd_sc_hd__inv_1
XFILLER_206_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$170 final_adder.U$$665/A final_adder.U$$664/A VGND VGND VPWR VPWR
+ final_adder.U$$276/A sky130_fd_sc_hd__and2_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$181 final_adder.U$$675/A final_adder.U$$547/B1 final_adder.U$$181/B1
+ VGND VGND VPWR VPWR final_adder.U$$181/X sky130_fd_sc_hd__a21o_1
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_1 dadda_fa_3_31_1/A dadda_fa_3_31_1/B dadda_fa_3_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_0/CIN dadda_fa_4_31_2/A sky130_fd_sc_hd__fa_1
XU$$3848 _554_/Q U$$3874/A2 U$$4259/B1 U$$3874/B2 VGND VGND VPWR VPWR U$$3849/A sky130_fd_sc_hd__a22o_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3859 U$$3859/A U$$3965/B VGND VGND VPWR VPWR U$$3859/X sky130_fd_sc_hd__xor2_1
XFILLER_206_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$192 final_adder.U$$687/A final_adder.U$$686/A VGND VGND VPWR VPWR
+ final_adder.U$$288/B sky130_fd_sc_hd__and2_1
XFILLER_205_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_24_0 U$$720/X U$$853/X U$$986/X VGND VGND VPWR VPWR dadda_fa_4_25_0/B
+ dadda_fa_4_24_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_526_ _526_/CLK _526_/D VGND VGND VPWR VPWR _526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_637 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_457_ _458_/CLK _457_/D VGND VGND VPWR VPWR _457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_388_ _520_/CLK _388_/D VGND VGND VPWR VPWR _388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_90_5 dadda_fa_2_90_5/A dadda_fa_2_90_5/B dadda_fa_2_90_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_91_2/A dadda_fa_4_90_0/A sky130_fd_sc_hd__fa_2
XFILLER_138_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_83_4 dadda_fa_2_83_4/A dadda_fa_2_83_4/B dadda_fa_2_83_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/CIN dadda_fa_3_83_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_76_3 dadda_fa_2_76_3/A dadda_fa_2_76_3/B dadda_fa_2_76_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/B dadda_fa_3_76_3/B sky130_fd_sc_hd__fa_1
XFILLER_130_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_69_2 dadda_fa_2_69_2/A dadda_fa_2_69_2/B dadda_fa_2_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/A dadda_fa_3_69_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_46_1 dadda_fa_5_46_1/A dadda_fa_5_46_1/B dadda_fa_5_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_47_0/B dadda_fa_7_46_0/A sky130_fd_sc_hd__fa_1
XFILLER_96_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_39_0 dadda_fa_5_39_0/A dadda_fa_5_39_0/B dadda_fa_5_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_40_0/A dadda_fa_6_39_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_37_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_120_1 dadda_fa_5_120_1/A dadda_fa_5_120_1/B dadda_ha_4_120_1/SUM VGND
+ VGND VPWR VPWR dadda_fa_6_121_0/B dadda_fa_7_120_0/A sky130_fd_sc_hd__fa_1
XFILLER_165_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_113_0 dadda_fa_5_113_0/A dadda_fa_5_113_0/B dadda_fa_5_113_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_114_0/A dadda_fa_6_113_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_71_2 U$$2942/X U$$3075/X U$$3208/X VGND VGND VPWR VPWR dadda_fa_2_72_1/A
+ dadda_fa_2_71_4/A sky130_fd_sc_hd__fa_1
XFILLER_28_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_64_1 U$$2928/X U$$3061/X U$$3194/X VGND VGND VPWR VPWR dadda_fa_2_65_0/CIN
+ dadda_fa_2_64_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_41_0 dadda_fa_4_41_0/A dadda_fa_4_41_0/B dadda_fa_4_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/A dadda_fa_5_41_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_57_0 U$$1185/X U$$1318/X U$$1451/X VGND VGND VPWR VPWR dadda_fa_2_58_0/B
+ dadda_fa_2_57_3/B sky130_fd_sc_hd__fa_1
XFILLER_46_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1709 U$$1709/A U$$1711/B VGND VGND VPWR VPWR U$$1709/X sky130_fd_sc_hd__xor2_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_311_ _444_/CLK _311_/D VGND VGND VPWR VPWR _311_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_242_ _372_/CLK _242_/D VGND VGND VPWR VPWR _242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1004 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_173_ _179_/CLK _173_/D VGND VGND VPWR VPWR _173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput19 a[26] VGND VGND VPWR VPWR _642_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_93_3 dadda_fa_3_93_3/A dadda_fa_3_93_3/B dadda_fa_3_93_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_1/B dadda_fa_4_93_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_328 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_86_2 dadda_fa_3_86_2/A dadda_fa_3_86_2/B dadda_fa_3_86_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_1/A dadda_fa_4_86_2/B sky130_fd_sc_hd__fa_1
XFILLER_123_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_79_1 dadda_fa_3_79_1/A dadda_fa_3_79_1/B dadda_fa_3_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_0/CIN dadda_fa_4_79_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_56_0 dadda_fa_6_56_0/A dadda_fa_6_56_0/B dadda_fa_6_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_57_0/B dadda_fa_7_56_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater609 U$$263/A2 VGND VGND VPWR VPWR U$$219/A2 sky130_fd_sc_hd__buf_6
XFILLER_42_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4302 U$$4302/A U$$4348/B VGND VGND VPWR VPWR U$$4302/X sky130_fd_sc_hd__xor2_1
XU$$4313 _581_/Q U$$4327/A2 _582_/Q U$$4333/B2 VGND VGND VPWR VPWR U$$4314/A sky130_fd_sc_hd__a22o_1
XFILLER_42_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4324 U$$4324/A U$$4334/B VGND VGND VPWR VPWR U$$4324/X sky130_fd_sc_hd__xor2_1
XFILLER_133_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4335 U$$4472/A1 U$$4335/A2 U$$4472/B1 U$$4252/X VGND VGND VPWR VPWR U$$4336/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3601 U$$3601/A U$$3637/B VGND VGND VPWR VPWR U$$3601/X sky130_fd_sc_hd__xor2_1
XU$$4346 U$$4346/A U$$4350/B VGND VGND VPWR VPWR U$$4346/X sky130_fd_sc_hd__xor2_1
XFILLER_203_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3612 U$$4160/A1 U$$3612/A2 U$$4160/B1 U$$3612/B2 VGND VGND VPWR VPWR U$$3613/A
+ sky130_fd_sc_hd__a22o_1
XU$$4357 U$$4357/A1 U$$4369/A2 U$$4494/B1 U$$4369/B2 VGND VGND VPWR VPWR U$$4358/A
+ sky130_fd_sc_hd__a22o_1
XU$$3623 U$$3623/A U$$3627/B VGND VGND VPWR VPWR U$$3623/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_115_2 dadda_fa_4_115_2/A dadda_fa_4_115_2/B dadda_fa_4_115_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_116_0/CIN dadda_fa_5_115_1/CIN sky130_fd_sc_hd__fa_1
XU$$4368 U$$4368/A U$$4384/A VGND VGND VPWR VPWR U$$4368/X sky130_fd_sc_hd__xor2_1
XU$$4379 U$$4516/A1 U$$4381/A2 U$$4516/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4380/A
+ sky130_fd_sc_hd__a22o_1
XU$$3634 U$$3769/B1 U$$3636/A2 U$$3771/B1 U$$3636/B2 VGND VGND VPWR VPWR U$$3635/A
+ sky130_fd_sc_hd__a22o_1
XU$$2900 U$$2900/A U$$2916/B VGND VGND VPWR VPWR U$$2900/X sky130_fd_sc_hd__xor2_1
XFILLER_19_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3645 U$$3645/A U$$3675/B VGND VGND VPWR VPWR U$$3645/X sky130_fd_sc_hd__xor2_1
XU$$3656 U$$3791/B1 U$$3664/A2 U$$3932/A1 U$$3664/B2 VGND VGND VPWR VPWR U$$3657/A
+ sky130_fd_sc_hd__a22o_1
XU$$2911 U$$3046/B1 U$$2981/A2 U$$310/A1 U$$2981/B2 VGND VGND VPWR VPWR U$$2912/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2922 U$$2922/A U$$2928/B VGND VGND VPWR VPWR U$$2922/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_108_1 dadda_fa_4_108_1/A dadda_fa_4_108_1/B dadda_fa_4_108_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/B dadda_fa_5_108_1/B sky130_fd_sc_hd__fa_1
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3667 U$$3667/A U$$3671/B VGND VGND VPWR VPWR U$$3667/X sky130_fd_sc_hd__xor2_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2933 U$$4301/B1 U$$2973/A2 U$$4305/A1 U$$2973/B2 VGND VGND VPWR VPWR U$$2934/A
+ sky130_fd_sc_hd__a22o_1
XU$$3678 U$$4361/B1 U$$3696/A2 U$$4502/A1 U$$3696/B2 VGND VGND VPWR VPWR U$$3679/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3689 U$$3689/A U$$3699/A VGND VGND VPWR VPWR U$$3689/X sky130_fd_sc_hd__xor2_1
XU$$2944 U$$2944/A U$$2944/B VGND VGND VPWR VPWR U$$2944/X sky130_fd_sc_hd__xor2_1
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2955 U$$4051/A1 U$$2997/A2 U$$2957/A1 U$$2997/B2 VGND VGND VPWR VPWR U$$2956/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2966 U$$2966/A U$$2966/B VGND VGND VPWR VPWR U$$2966/X sky130_fd_sc_hd__xor2_1
XFILLER_206_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2977 U$$922/A1 U$$2981/A2 U$$3799/B1 U$$2981/B2 VGND VGND VPWR VPWR U$$2978/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_260 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_271 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2988 U$$2988/A U$$2988/B VGND VGND VPWR VPWR U$$2988/X sky130_fd_sc_hd__xor2_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_509_ _510_/CLK _509_/D VGND VGND VPWR VPWR _509_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2999 _609_/Q U$$3005/A2 U$$2999/B1 U$$3005/B2 VGND VGND VPWR VPWR U$$3000/A sky130_fd_sc_hd__a22o_1
XANTENNA_282 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_293 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_81_1 dadda_fa_2_81_1/A dadda_fa_2_81_1/B dadda_fa_2_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_0/CIN dadda_fa_3_81_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_74_0 dadda_fa_2_74_0/A dadda_fa_2_74_0/B dadda_fa_2_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_0/B dadda_fa_3_74_2/B sky130_fd_sc_hd__fa_1
XFILLER_114_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_50_7 U$$2900/X U$$3033/X U$$3166/X VGND VGND VPWR VPWR dadda_fa_2_51_2/CIN
+ dadda_fa_2_50_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_96_1 dadda_fa_4_96_1/A dadda_fa_4_96_1/B dadda_fa_4_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/B dadda_fa_5_96_1/B sky130_fd_sc_hd__fa_1
XFILLER_125_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_73_0 dadda_fa_7_73_0/A dadda_fa_7_73_0/B dadda_fa_7_73_0/CIN VGND VGND
+ VPWR VPWR _498_/D _369_/D sky130_fd_sc_hd__fa_1
XFILLER_156_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_89_0 dadda_fa_4_89_0/A dadda_fa_4_89_0/B dadda_fa_4_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/A dadda_fa_5_89_1/A sky130_fd_sc_hd__fa_1
XFILLER_152_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2207 U$$2207/A U$$2241/B VGND VGND VPWR VPWR U$$2207/X sky130_fd_sc_hd__xor2_1
XFILLER_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2218 U$$3451/A1 U$$2262/A2 U$$3453/A1 U$$2262/B2 VGND VGND VPWR VPWR U$$2219/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_784 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2229 U$$2229/A U$$2243/B VGND VGND VPWR VPWR U$$2229/X sky130_fd_sc_hd__xor2_1
XFILLER_15_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1506 U$$1507/A VGND VGND VPWR VPWR U$$1506/Y sky130_fd_sc_hd__inv_1
XFILLER_167_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1517 U$$695/A1 U$$1557/A2 U$$2613/B1 U$$1557/B2 VGND VGND VPWR VPWR U$$1518/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_1134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1528 U$$1528/A U$$1554/B VGND VGND VPWR VPWR U$$1528/X sky130_fd_sc_hd__xor2_1
XFILLER_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1539 U$$2909/A1 U$$1577/A2 U$$2909/B1 U$$1577/B2 VGND VGND VPWR VPWR U$$1540/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_467 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_225_ _225_/CLK _225_/D VGND VGND VPWR VPWR _225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_91_0 dadda_fa_3_91_0/A dadda_fa_3_91_0/B dadda_fa_3_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_0/B dadda_fa_4_91_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater406 U$$795/A2 VGND VGND VPWR VPWR U$$759/A2 sky130_fd_sc_hd__buf_6
Xrepeater417 U$$4251/X VGND VGND VPWR VPWR U$$4297/A2 sky130_fd_sc_hd__buf_6
Xrepeater428 U$$415/X VGND VGND VPWR VPWR U$$491/A2 sky130_fd_sc_hd__buf_4
XU$$4110 _675_/Q VGND VGND VPWR VPWR U$$4110/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_2_53_5 dadda_fa_2_53_5/A dadda_fa_2_53_5/B dadda_fa_2_53_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_2/A dadda_fa_4_53_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_120_0 dadda_fa_4_120_0/A U$$3971/X U$$4104/X VGND VGND VPWR VPWR dadda_fa_5_121_1/A
+ dadda_fa_5_120_1/B sky130_fd_sc_hd__fa_1
XFILLER_93_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater439 U$$52/A2 VGND VGND VPWR VPWR U$$8/A2 sky130_fd_sc_hd__clkbuf_4
XU$$4121 U$$4121/A U$$4141/B VGND VGND VPWR VPWR U$$4121/X sky130_fd_sc_hd__xor2_1
XU$$4132 U$$4269/A1 U$$4226/A2 _560_/Q U$$4226/B2 VGND VGND VPWR VPWR U$$4133/A sky130_fd_sc_hd__a22o_1
XU$$4143 U$$4143/A U$$4183/B VGND VGND VPWR VPWR U$$4143/X sky130_fd_sc_hd__xor2_1
XU$$4154 U$$4154/A1 U$$4182/A2 U$$4154/B1 U$$4182/B2 VGND VGND VPWR VPWR U$$4155/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3420 U$$4516/A1 U$$3292/X U$$4516/B1 U$$3293/X VGND VGND VPWR VPWR U$$3421/A sky130_fd_sc_hd__a22o_1
XU$$4165 U$$4165/A U$$4175/B VGND VGND VPWR VPWR U$$4165/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_46_4 dadda_fa_2_46_4/A dadda_fa_2_46_4/B dadda_fa_2_46_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/CIN dadda_fa_3_46_3/CIN sky130_fd_sc_hd__fa_1
XU$$3431 U$$3431/A1 U$$3479/A2 U$$3844/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3432/A
+ sky130_fd_sc_hd__a22o_1
XU$$4176 U$$4176/A1 U$$4202/A2 U$$4176/B1 U$$4202/B2 VGND VGND VPWR VPWR U$$4177/A
+ sky130_fd_sc_hd__a22o_1
XU$$4187 U$$4187/A U$$4197/B VGND VGND VPWR VPWR U$$4187/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3442 U$$3442/A U$$3490/B VGND VGND VPWR VPWR U$$3442/X sky130_fd_sc_hd__xor2_1
XFILLER_25_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4198 U$$4333/B1 U$$4202/A2 U$$4198/B1 U$$4202/B2 VGND VGND VPWR VPWR U$$4199/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3453 U$$3453/A1 U$$3497/A2 U$$3453/B1 U$$3497/B2 VGND VGND VPWR VPWR U$$3454/A
+ sky130_fd_sc_hd__a22o_1
XU$$3464 U$$3464/A U$$3561/A VGND VGND VPWR VPWR U$$3464/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_39_3 U$$2346/X U$$2479/X U$$2612/X VGND VGND VPWR VPWR dadda_fa_3_40_1/B
+ dadda_fa_3_39_3/B sky130_fd_sc_hd__fa_1
XU$$2730 U$$2730/A U$$2730/B VGND VGND VPWR VPWR U$$2730/X sky130_fd_sc_hd__xor2_1
XU$$3475 U$$3475/A1 U$$3479/A2 U$$3475/B1 U$$3479/B2 VGND VGND VPWR VPWR U$$3476/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2741 _656_/Q VGND VGND VPWR VPWR U$$2743/B sky130_fd_sc_hd__inv_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3486 U$$3486/A U$$3490/B VGND VGND VPWR VPWR U$$3486/X sky130_fd_sc_hd__xor2_1
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2752 U$$3024/B1 U$$2798/A2 U$$2754/A1 U$$2798/B2 VGND VGND VPWR VPWR U$$2753/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3497 U$$4045/A1 U$$3497/A2 U$$4456/B1 U$$3497/B2 VGND VGND VPWR VPWR U$$3498/A
+ sky130_fd_sc_hd__a22o_1
XU$$2763 U$$2763/A U$$2813/B VGND VGND VPWR VPWR U$$2763/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2774 U$$2909/B1 U$$2814/A2 U$$2774/B1 U$$2814/B2 VGND VGND VPWR VPWR U$$2775/A
+ sky130_fd_sc_hd__a22o_1
XU$$2785 U$$2785/A U$$2787/B VGND VGND VPWR VPWR U$$2785/X sky130_fd_sc_hd__xor2_1
XU$$2796 U$$4301/B1 U$$2798/A2 U$$2796/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2797/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_976 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput209 c[57] VGND VGND VPWR VPWR input209/X sky130_fd_sc_hd__clkbuf_4
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$703 final_adder.U$$703/A final_adder.U$$703/B VGND VGND VPWR VPWR
+ _249_/D sky130_fd_sc_hd__xor2_1
XTAP_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$714 final_adder.U$$714/A final_adder.U$$714/B VGND VGND VPWR VPWR
+ _260_/D sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$725 final_adder.U$$725/A final_adder.U$$725/B VGND VGND VPWR VPWR
+ _271_/D sky130_fd_sc_hd__xor2_1
XFILLER_151_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$736 final_adder.U$$736/A final_adder.U$$736/B VGND VGND VPWR VPWR
+ _282_/D sky130_fd_sc_hd__xor2_4
XFILLER_84_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater940 U$$3764/B VGND VGND VPWR VPWR U$$3760/B sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$747 final_adder.U$$747/A final_adder.U$$747/B VGND VGND VPWR VPWR
+ _293_/D sky130_fd_sc_hd__xor2_4
Xrepeater951 _669_/Q VGND VGND VPWR VPWR U$$3698/A sky130_fd_sc_hd__buf_6
XFILLER_83_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater962 U$$3520/B VGND VGND VPWR VPWR U$$3490/B sky130_fd_sc_hd__buf_6
XU$$608 U$$745/A1 U$$616/A2 U$$882/B1 U$$616/B2 VGND VGND VPWR VPWR U$$609/A sky130_fd_sc_hd__a22o_1
Xrepeater973 U$$3425/A VGND VGND VPWR VPWR U$$3407/B sky130_fd_sc_hd__buf_6
XFILLER_99_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$619 U$$619/A U$$669/B VGND VGND VPWR VPWR U$$619/X sky130_fd_sc_hd__xor2_1
Xrepeater984 U$$3107/B VGND VGND VPWR VPWR U$$3065/B sky130_fd_sc_hd__buf_6
XFILLER_95_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater995 U$$2982/B VGND VGND VPWR VPWR U$$2988/B sky130_fd_sc_hd__buf_6
XFILLER_17_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_47 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1508 _576_/Q VGND VGND VPWR VPWR U$$3618/A1 sky130_fd_sc_hd__buf_4
XFILLER_116_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1519 U$$3342/A1 VGND VGND VPWR VPWR U$$52/B1 sky130_fd_sc_hd__buf_6
XFILLER_119_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_108_0 U$$3282/X U$$3415/X U$$3548/X VGND VGND VPWR VPWR dadda_fa_4_109_0/B
+ dadda_fa_4_108_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_56_3 dadda_fa_3_56_3/A dadda_fa_3_56_3/B dadda_fa_3_56_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_1/B dadda_fa_4_56_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_616 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_49_2 dadda_fa_3_49_2/A dadda_fa_3_49_2/B dadda_fa_3_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_1/A dadda_fa_4_49_2/B sky130_fd_sc_hd__fa_1
XFILLER_208_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2004 U$$3783/B1 U$$2040/A2 U$$2963/B1 U$$2040/B2 VGND VGND VPWR VPWR U$$2005/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2015 U$$2015/A U$$2029/B VGND VGND VPWR VPWR U$$2015/X sky130_fd_sc_hd__xor2_1
XFILLER_207_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2026 U$$3122/A1 U$$2052/A2 U$$382/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2027/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_19_0 dadda_fa_6_19_0/A dadda_fa_6_19_0/B dadda_fa_6_19_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_20_0/B dadda_fa_7_19_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_74_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2037 U$$2037/A U$$2039/B VGND VGND VPWR VPWR U$$2037/X sky130_fd_sc_hd__xor2_1
XU$$1303 U$$344/A1 U$$1309/A2 U$$72/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1304/A sky130_fd_sc_hd__a22o_1
XU$$2048 U$$3418/A1 U$$2052/A2 U$$2459/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2049/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1314 U$$1314/A U$$1356/B VGND VGND VPWR VPWR U$$1314/X sky130_fd_sc_hd__xor2_1
XU$$2059 U$$2057/Y _646_/Q _645_/Q U$$2058/X U$$2055/Y VGND VGND VPWR VPWR U$$2059/X
+ sky130_fd_sc_hd__a32o_4
XU$$1325 U$$92/A1 U$$1237/X U$$94/A1 U$$1238/X VGND VGND VPWR VPWR U$$1326/A sky130_fd_sc_hd__a22o_1
XU$$1336 U$$1336/A U$$1370/A VGND VGND VPWR VPWR U$$1336/X sky130_fd_sc_hd__xor2_1
XU$$1347 U$$251/A1 U$$1355/A2 U$$251/B1 U$$1355/B2 VGND VGND VPWR VPWR U$$1348/A sky130_fd_sc_hd__a22o_1
XFILLER_16_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1358 U$$1358/A U$$1368/B VGND VGND VPWR VPWR U$$1358/X sky130_fd_sc_hd__xor2_1
XFILLER_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1369 U$$1369/A VGND VGND VPWR VPWR U$$1369/Y sky130_fd_sc_hd__inv_1
XFILLER_128_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_208_ _478_/CLK _208_/D VGND VGND VPWR VPWR _208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_718 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_51_2 dadda_fa_2_51_2/A dadda_fa_2_51_2/B dadda_fa_2_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/A dadda_fa_3_51_3/A sky130_fd_sc_hd__fa_1
XFILLER_22_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_44_1 U$$2755/X U$$2888/X U$$3021/X VGND VGND VPWR VPWR dadda_fa_3_45_0/CIN
+ dadda_fa_3_44_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$10 _434_/Q _306_/Q VGND VGND VPWR VPWR final_adder.U$$505/B1 final_adder.U$$632/A
+ sky130_fd_sc_hd__ha_2
XU$$3250 U$$3250/A U$$3256/B VGND VGND VPWR VPWR U$$3250/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$21 _445_/Q _317_/Q VGND VGND VPWR VPWR final_adder.U$$149/B1 final_adder.U$$643/A
+ sky130_fd_sc_hd__ha_2
Xdadda_fa_5_21_0 dadda_fa_5_21_0/A dadda_fa_5_21_0/B dadda_fa_5_21_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_22_0/A dadda_fa_6_21_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$32 _456_/Q _328_/Q VGND VGND VPWR VPWR final_adder.U$$527/B1 final_adder.U$$654/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_2_37_0 U$$746/X U$$879/X U$$1012/X VGND VGND VPWR VPWR dadda_fa_3_38_0/B
+ dadda_fa_3_37_2/B sky130_fd_sc_hd__fa_1
XU$$3261 _603_/Q U$$3263/A2 _604_/Q U$$3263/B2 VGND VGND VPWR VPWR U$$3262/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$43 _467_/Q _339_/Q VGND VGND VPWR VPWR final_adder.U$$171/B1 final_adder.U$$665/A
+ sky130_fd_sc_hd__ha_1
XFILLER_53_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3272 U$$3272/A U$$3272/B VGND VGND VPWR VPWR U$$3272/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$54 _478_/Q _350_/Q VGND VGND VPWR VPWR final_adder.U$$549/B1 final_adder.U$$676/A
+ sky130_fd_sc_hd__ha_1
XU$$3283 U$$3283/A1 U$$3283/A2 U$$3285/A1 U$$3283/B2 VGND VGND VPWR VPWR U$$3284/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$65 _489_/Q _361_/Q VGND VGND VPWR VPWR final_adder.U$$193/B1 final_adder.U$$687/A
+ sky130_fd_sc_hd__ha_2
XU$$3294 U$$3294/A1 U$$3320/A2 _552_/Q U$$3320/B2 VGND VGND VPWR VPWR U$$3295/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$76 _500_/Q _372_/Q VGND VGND VPWR VPWR final_adder.U$$571/B1 final_adder.U$$698/A
+ sky130_fd_sc_hd__ha_1
XU$$2560 U$$916/A1 U$$2566/A2 U$$3519/B1 U$$2566/B2 VGND VGND VPWR VPWR U$$2561/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$87 _511_/Q _383_/Q VGND VGND VPWR VPWR final_adder.U$$215/B1 final_adder.U$$709/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$98 _522_/Q _394_/Q VGND VGND VPWR VPWR final_adder.U$$593/B1 final_adder.U$$720/A
+ sky130_fd_sc_hd__ha_1
XFILLER_146_1132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2571 U$$2571/A _653_/Q VGND VGND VPWR VPWR U$$2571/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2582 U$$3404/A1 U$$2600/A2 U$$3132/A1 U$$2600/B2 VGND VGND VPWR VPWR U$$2583/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2593 U$$2593/A U$$2597/B VGND VGND VPWR VPWR U$$2593/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1870 U$$1870/A U$$1870/B VGND VGND VPWR VPWR U$$1870/X sky130_fd_sc_hd__xor2_1
XFILLER_179_578 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1881 U$$98/B1 U$$1915/A2 U$$785/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1882/A sky130_fd_sc_hd__a22o_1
XU$$1892 U$$1892/A U$$1917/A VGND VGND VPWR VPWR U$$1892/X sky130_fd_sc_hd__xor2_1
XFILLER_142_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$554_1840 VGND VGND VPWR VPWR U$$554_1840/HI U$$554/A1 sky130_fd_sc_hd__conb_1
XFILLER_116_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_810 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_89_3 U$$2978/X U$$3111/X U$$3244/X VGND VGND VPWR VPWR dadda_fa_2_90_4/CIN
+ dadda_fa_3_89_0/A sky130_fd_sc_hd__fa_1
XFILLER_153_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_66_2 dadda_fa_4_66_2/A dadda_fa_4_66_2/B dadda_fa_4_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/CIN dadda_fa_5_66_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_59_1 dadda_fa_4_59_1/A dadda_fa_4_59_1/B dadda_fa_4_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/B dadda_fa_5_59_1/B sky130_fd_sc_hd__fa_1
XTAP_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_36_0 dadda_fa_7_36_0/A dadda_fa_7_36_0/B dadda_fa_7_36_0/CIN VGND VGND
+ VPWR VPWR _461_/D _332_/D sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$511 final_adder.U$$638/A final_adder.U$$638/B final_adder.U$$511/B1
+ VGND VGND VPWR VPWR final_adder.U$$639/B sky130_fd_sc_hd__a21o_1
XTAP_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$533 final_adder.U$$660/A final_adder.U$$660/B final_adder.U$$533/B1
+ VGND VGND VPWR VPWR final_adder.U$$661/B sky130_fd_sc_hd__a21o_1
XTAP_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$555 final_adder.U$$682/A final_adder.U$$682/B final_adder.U$$555/B1
+ VGND VGND VPWR VPWR final_adder.U$$683/B sky130_fd_sc_hd__a21o_1
XFILLER_151_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$405 U$$405/A U$$411/A VGND VGND VPWR VPWR U$$405/X sky130_fd_sc_hd__xor2_1
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater770 U$$408/B2 VGND VGND VPWR VPWR U$$398/B2 sky130_fd_sc_hd__buf_4
XFILLER_45_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$577 final_adder.U$$704/A final_adder.U$$704/B final_adder.U$$577/B1
+ VGND VGND VPWR VPWR final_adder.U$$705/B sky130_fd_sc_hd__a21o_1
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$416 U$$414/B U$$411/A _622_/Q U$$411/Y VGND VGND VPWR VPWR U$$416/X sky130_fd_sc_hd__a22o_4
XFILLER_56_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater781 U$$2874/B2 VGND VGND VPWR VPWR U$$2866/B2 sky130_fd_sc_hd__clkbuf_8
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$427 U$$973/B1 U$$447/A2 U$$429/A1 U$$447/B2 VGND VGND VPWR VPWR U$$428/A sky130_fd_sc_hd__a22o_1
Xrepeater792 U$$2471/X VGND VGND VPWR VPWR U$$2566/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$599 final_adder.U$$726/A final_adder.U$$726/B final_adder.U$$599/B1
+ VGND VGND VPWR VPWR final_adder.U$$727/B sky130_fd_sc_hd__a21o_1
XU$$438 U$$438/A U$$456/B VGND VGND VPWR VPWR U$$438/X sky130_fd_sc_hd__xor2_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$449 U$$449/A1 U$$483/A2 U$$449/B1 U$$483/B2 VGND VGND VPWR VPWR U$$450/A sky130_fd_sc_hd__a22o_1
X_490_ _491_/CLK _490_/D VGND VGND VPWR VPWR _490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1305 _602_/Q VGND VGND VPWR VPWR U$$3805/B1 sky130_fd_sc_hd__buf_6
XFILLER_165_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1316 U$$3253/B1 VGND VGND VPWR VPWR U$$2431/B1 sky130_fd_sc_hd__buf_6
XFILLER_138_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1327 _599_/Q VGND VGND VPWR VPWR U$$3799/B1 sky130_fd_sc_hd__buf_4
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1338 _598_/Q VGND VGND VPWR VPWR U$$3934/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_153_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1349 U$$3932/A1 VGND VGND VPWR VPWR U$$96/A1 sky130_fd_sc_hd__buf_4
XFILLER_119_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_61_1 dadda_fa_3_61_1/A dadda_fa_3_61_1/B dadda_fa_3_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_0/CIN dadda_fa_4_61_2/A sky130_fd_sc_hd__fa_1
XFILLER_192_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_54_0 dadda_fa_3_54_0/A dadda_fa_3_54_0/B dadda_fa_3_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_0/B dadda_fa_4_54_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_443 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$950 U$$950/A1 U$$956/A2 U$$950/B1 U$$956/B2 VGND VGND VPWR VPWR U$$951/A sky130_fd_sc_hd__a22o_1
XFILLER_211_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1100 U$$1098/Y _632_/Q _631_/Q U$$1099/X U$$1096/Y VGND VGND VPWR VPWR U$$1100/X
+ sky130_fd_sc_hd__a32o_1
XU$$961 _631_/Q VGND VGND VPWR VPWR U$$961/Y sky130_fd_sc_hd__inv_1
XFILLER_141_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1111 U$$1111/A U$$1147/B VGND VGND VPWR VPWR U$$1111/X sky130_fd_sc_hd__xor2_1
XU$$972 U$$972/A U$$994/B VGND VGND VPWR VPWR U$$972/X sky130_fd_sc_hd__xor2_1
XU$$1122 U$$985/A1 U$$1150/A2 U$$987/A1 U$$1150/B2 VGND VGND VPWR VPWR U$$1123/A sky130_fd_sc_hd__a22o_1
XU$$983 U$$24/A1 U$$997/A2 U$$985/A1 U$$997/B2 VGND VGND VPWR VPWR U$$984/A sky130_fd_sc_hd__a22o_1
XU$$994 U$$994/A U$$994/B VGND VGND VPWR VPWR U$$994/X sky130_fd_sc_hd__xor2_1
XU$$1133 U$$1133/A U$$1151/B VGND VGND VPWR VPWR U$$1133/X sky130_fd_sc_hd__xor2_1
XU$$1144 U$$48/A1 U$$1146/A2 U$$48/B1 U$$1146/B2 VGND VGND VPWR VPWR U$$1145/A sky130_fd_sc_hd__a22o_1
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1155 U$$1155/A U$$1195/B VGND VGND VPWR VPWR U$$1155/X sky130_fd_sc_hd__xor2_1
XFILLER_189_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1166 U$$3358/A1 U$$1176/A2 U$$894/A1 U$$1176/B2 VGND VGND VPWR VPWR U$$1167/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1177 U$$1177/A U$$1177/B VGND VGND VPWR VPWR U$$1177/X sky130_fd_sc_hd__xor2_1
XFILLER_149_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1188 U$$229/A1 U$$1208/A2 U$$2832/B1 U$$1208/B2 VGND VGND VPWR VPWR U$$1189/A
+ sky130_fd_sc_hd__a22o_1
XU$$1199 U$$1199/A U$$1203/B VGND VGND VPWR VPWR U$$1199/X sky130_fd_sc_hd__xor2_1
XFILLER_148_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_111_0 dadda_fa_7_111_0/A dadda_fa_7_111_0/B dadda_fa_7_111_0/CIN VGND
+ VGND VPWR VPWR _536_/D _407_/D sky130_fd_sc_hd__fa_1
XFILLER_54_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_99_2 U$$3264/X U$$3397/X U$$3530/X VGND VGND VPWR VPWR dadda_fa_3_100_1/CIN
+ dadda_fa_3_99_3/B sky130_fd_sc_hd__fa_1
Xdadda_fa_5_76_1 dadda_fa_5_76_1/A dadda_fa_5_76_1/B dadda_fa_5_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_77_0/B dadda_fa_7_76_0/A sky130_fd_sc_hd__fa_1
XFILLER_104_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_692 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_69_0 dadda_fa_5_69_0/A dadda_fa_5_69_0/B dadda_fa_5_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_70_0/A dadda_fa_6_69_0/CIN sky130_fd_sc_hd__fa_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_8 dadda_fa_1_68_8/A dadda_fa_1_68_8/B dadda_fa_1_68_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_3/A dadda_fa_3_68_0/A sky130_fd_sc_hd__fa_1
XFILLER_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$545_1839 VGND VGND VPWR VPWR U$$545_1839/HI U$$545/B1 sky130_fd_sc_hd__conb_1
XU$$3080 U$$3217/A1 U$$3082/A2 U$$4450/B1 U$$3082/B2 VGND VGND VPWR VPWR U$$3081/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3091 U$$3091/A U$$3111/B VGND VGND VPWR VPWR U$$3091/X sky130_fd_sc_hd__xor2_1
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_8_0 dadda_fa_6_8_0/A dadda_fa_6_8_0/B dadda_fa_6_8_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_9_0/B dadda_fa_7_8_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_198_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2390 U$$2390/A U$$2400/B VGND VGND VPWR VPWR U$$2390/X sky130_fd_sc_hd__xor2_1
XFILLER_10_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_71_0 dadda_fa_4_71_0/A dadda_fa_4_71_0/B dadda_fa_4_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/A dadda_fa_5_71_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_87_0 U$$1643/Y U$$1777/X U$$1910/X VGND VGND VPWR VPWR dadda_fa_2_88_3/A
+ dadda_fa_2_87_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1019 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$330 final_adder.U$$330/A final_adder.U$$330/B VGND VGND VPWR VPWR
+ final_adder.U$$356/A sky130_fd_sc_hd__and2_1
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_611_ _615_/CLK _611_/D VGND VGND VPWR VPWR _611_/Q sky130_fd_sc_hd__dfxtp_4
Xfinal_adder.U$$341 final_adder.U$$340/A final_adder.U$$297/X final_adder.U$$299/X
+ VGND VGND VPWR VPWR final_adder.U$$341/X sky130_fd_sc_hd__a21o_1
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_922 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$363 final_adder.U$$362/A final_adder.U$$341/X final_adder.U$$343/X
+ VGND VGND VPWR VPWR final_adder.U$$363/X sky130_fd_sc_hd__a21o_1
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$202 U$$202/A U$$232/B VGND VGND VPWR VPWR U$$202/X sky130_fd_sc_hd__xor2_1
XU$$213 U$$76/A1 U$$217/A2 U$$78/A1 U$$217/B2 VGND VGND VPWR VPWR U$$214/A sky130_fd_sc_hd__a22o_1
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$385 final_adder.U$$370/B final_adder.U$$654/B final_adder.U$$357/X
+ VGND VGND VPWR VPWR final_adder.U$$670/B sky130_fd_sc_hd__a21o_1
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$224 U$$224/A U$$226/B VGND VGND VPWR VPWR U$$224/X sky130_fd_sc_hd__xor2_1
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_542_ _542_/CLK _542_/D VGND VGND VPWR VPWR _542_/Q sky130_fd_sc_hd__dfxtp_1
XU$$235 U$$98/A1 U$$249/A2 U$$98/B1 U$$249/B2 VGND VGND VPWR VPWR U$$236/A sky130_fd_sc_hd__a22o_1
XU$$246 U$$246/A U$$250/B VGND VGND VPWR VPWR U$$246/X sky130_fd_sc_hd__xor2_1
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$257 U$$942/A1 U$$259/A2 U$$942/B1 U$$259/B2 VGND VGND VPWR VPWR U$$258/A sky130_fd_sc_hd__a22o_1
XFILLER_73_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$268 U$$268/A U$$272/B VGND VGND VPWR VPWR U$$268/X sky130_fd_sc_hd__xor2_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$279 U$$277/B _619_/Q _620_/Q U$$274/Y VGND VGND VPWR VPWR U$$279/X sky130_fd_sc_hd__a22o_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_473_ _475_/CLK _473_/D VGND VGND VPWR VPWR _473_/Q sky130_fd_sc_hd__dfxtp_1
XU$$4505_1831 VGND VGND VPWR VPWR U$$4505_1831/HI U$$4505/B sky130_fd_sc_hd__conb_1
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_75 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$7 U$$7/A U$$9/B VGND VGND VPWR VPWR U$$7/X sky130_fd_sc_hd__xor2_1
XFILLER_5_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_86_0 dadda_fa_6_86_0/A dadda_fa_6_86_0/B dadda_fa_6_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_87_0/B dadda_fa_7_86_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1102 U$$1369/A VGND VGND VPWR VPWR U$$1368/B sky130_fd_sc_hd__buf_8
Xrepeater1113 U$$1191/B VGND VGND VPWR VPWR U$$1177/B sky130_fd_sc_hd__buf_6
XFILLER_154_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1124 U$$998/B VGND VGND VPWR VPWR U$$982/B sky130_fd_sc_hd__buf_6
XFILLER_126_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1135 U$$951/B VGND VGND VPWR VPWR U$$958/A sky130_fd_sc_hd__buf_6
XFILLER_153_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1146 _627_/Q VGND VGND VPWR VPWR U$$804/B sky130_fd_sc_hd__buf_6
Xrepeater1157 U$$500/B VGND VGND VPWR VPWR U$$452/B sky130_fd_sc_hd__buf_6
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1168 U$$383/B VGND VGND VPWR VPWR U$$351/B sky130_fd_sc_hd__buf_12
Xrepeater1179 U$$264/B VGND VGND VPWR VPWR U$$232/B sky130_fd_sc_hd__buf_12
XFILLER_153_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_662 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$780 U$$780/A U$$816/B VGND VGND VPWR VPWR U$$780/X sky130_fd_sc_hd__xor2_1
XFILLER_211_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$791 U$$791/A1 U$$809/A2 U$$791/B1 U$$809/B2 VGND VGND VPWR VPWR U$$792/A sky130_fd_sc_hd__a22o_1
XFILLER_108_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_80_7 U$$3891/X U$$4024/X U$$4157/X VGND VGND VPWR VPWR dadda_fa_2_81_3/A
+ dadda_fa_2_80_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1680 U$$3163/B1 VGND VGND VPWR VPWR U$$2343/A1 sky130_fd_sc_hd__buf_4
XFILLER_28_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1691 U$$2478/A1 VGND VGND VPWR VPWR U$$12/A1 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_1_73_6 U$$4276/X U$$4409/X input227/X VGND VGND VPWR VPWR dadda_fa_2_74_2/B
+ dadda_fa_2_73_5/B sky130_fd_sc_hd__fa_1
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_66_5 input219/X dadda_fa_1_66_5/B dadda_fa_1_66_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_67_2/A dadda_fa_2_66_5/A sky130_fd_sc_hd__fa_2
XFILLER_86_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_59_4 U$$3184/X U$$3317/X U$$3450/X VGND VGND VPWR VPWR dadda_fa_2_60_1/CIN
+ dadda_fa_2_59_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_443 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_29_2 dadda_fa_4_29_2/A dadda_fa_4_29_2/B dadda_fa_4_29_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/CIN dadda_fa_5_29_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_187_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_805 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4506 U$$4506/A1 U$$4388/X U$$4508/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4507/A
+ sky130_fd_sc_hd__a22o_1
XU$$4517 U$$4517/A U$$4517/B VGND VGND VPWR VPWR U$$4517/X sky130_fd_sc_hd__xor2_1
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3805 U$$3805/A1 U$$3805/A2 U$$3805/B1 U$$3805/B2 VGND VGND VPWR VPWR U$$3806/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_3_18_2 U$$841/X U$$974/X VGND VGND VPWR VPWR dadda_fa_4_19_1/CIN dadda_ha_3_18_2/SUM
+ sky130_fd_sc_hd__ha_1
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3816 U$$3816/A U$$3816/B VGND VGND VPWR VPWR U$$3816/X sky130_fd_sc_hd__xor2_1
XFILLER_64_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3827 U$$4238/A1 U$$3833/A2 U$$4238/B1 U$$3833/B2 VGND VGND VPWR VPWR U$$3828/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$160 final_adder.U$$655/A final_adder.U$$654/A VGND VGND VPWR VPWR
+ final_adder.U$$272/B sky130_fd_sc_hd__and2_1
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3838 _673_/Q VGND VGND VPWR VPWR U$$3838/Y sky130_fd_sc_hd__inv_1
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$171 final_adder.U$$665/A final_adder.U$$537/B1 final_adder.U$$171/B1
+ VGND VGND VPWR VPWR final_adder.U$$171/X sky130_fd_sc_hd__a21o_1
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3849 U$$3849/A U$$3873/B VGND VGND VPWR VPWR U$$3849/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$182 final_adder.U$$677/A final_adder.U$$676/A VGND VGND VPWR VPWR
+ final_adder.U$$282/A sky130_fd_sc_hd__and2_1
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_31_2 dadda_fa_3_31_2/A dadda_fa_3_31_2/B dadda_fa_3_31_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_1/A dadda_fa_4_31_2/B sky130_fd_sc_hd__fa_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$193 final_adder.U$$687/A final_adder.U$$559/B1 final_adder.U$$193/B1
+ VGND VGND VPWR VPWR final_adder.U$$193/X sky130_fd_sc_hd__a21o_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_24_1 U$$1119/X U$$1252/X U$$1385/X VGND VGND VPWR VPWR dadda_fa_4_25_0/CIN
+ dadda_fa_4_24_2/A sky130_fd_sc_hd__fa_1
XFILLER_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_525_ _535_/CLK _525_/D VGND VGND VPWR VPWR _525_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_17_0 U$$41/X U$$174/X U$$307/X VGND VGND VPWR VPWR dadda_fa_4_18_1/B dadda_fa_4_17_2/B
+ sky130_fd_sc_hd__fa_1
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_456_ _478_/CLK _456_/D VGND VGND VPWR VPWR _456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_387_ _560_/CLK _387_/D VGND VGND VPWR VPWR _387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_83_5 dadda_fa_2_83_5/A dadda_fa_2_83_5/B dadda_fa_2_83_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_2/A dadda_fa_4_83_0/A sky130_fd_sc_hd__fa_2
XFILLER_114_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_76_4 dadda_fa_2_76_4/A dadda_fa_2_76_4/B dadda_fa_2_76_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/CIN dadda_fa_3_76_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_971 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_69_3 dadda_fa_2_69_3/A dadda_fa_2_69_3/B dadda_fa_2_69_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/B dadda_fa_3_69_3/B sky130_fd_sc_hd__fa_1
XFILLER_110_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_39_1 dadda_fa_5_39_1/A dadda_fa_5_39_1/B dadda_fa_5_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_40_0/B dadda_fa_7_39_0/A sky130_fd_sc_hd__fa_2
XFILLER_23_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_113_1 dadda_fa_5_113_1/A dadda_fa_5_113_1/B dadda_fa_5_113_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_114_0/B dadda_fa_7_113_0/A sky130_fd_sc_hd__fa_1
XFILLER_176_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_106_0 dadda_fa_5_106_0/A dadda_fa_5_106_0/B dadda_fa_5_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_107_0/A dadda_fa_6_106_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_71_3 U$$3341/X U$$3474/X U$$3607/X VGND VGND VPWR VPWR dadda_fa_2_72_1/B
+ dadda_fa_2_71_4/B sky130_fd_sc_hd__fa_1
XFILLER_113_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_64_2 U$$3327/X U$$3460/X U$$3593/X VGND VGND VPWR VPWR dadda_fa_2_65_1/A
+ dadda_fa_2_64_4/A sky130_fd_sc_hd__fa_1
XFILLER_59_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_41_1 dadda_fa_4_41_1/A dadda_fa_4_41_1/B dadda_fa_4_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/B dadda_fa_5_41_1/B sky130_fd_sc_hd__fa_1
XFILLER_28_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_57_1 U$$1584/X U$$1717/X U$$1850/X VGND VGND VPWR VPWR dadda_fa_2_58_0/CIN
+ dadda_fa_2_57_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_34_0 dadda_fa_4_34_0/A dadda_fa_4_34_0/B dadda_fa_4_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/A dadda_fa_5_34_1/A sky130_fd_sc_hd__fa_1
XFILLER_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_310_ _439_/CLK _310_/D VGND VGND VPWR VPWR _310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_241_ _503_/CLK _241_/D VGND VGND VPWR VPWR _241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_172_ _179_/CLK _172_/D VGND VGND VPWR VPWR _172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_86_3 dadda_fa_3_86_3/A dadda_fa_3_86_3/B dadda_fa_3_86_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_1/B dadda_fa_4_86_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_184_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_79_2 dadda_fa_3_79_2/A dadda_fa_3_79_2/B dadda_fa_3_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_1/A dadda_fa_4_79_2/B sky130_fd_sc_hd__fa_1
XFILLER_112_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_49_0 dadda_fa_6_49_0/A dadda_fa_6_49_0/B dadda_fa_6_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_50_0/B dadda_fa_7_49_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_38_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4303 U$$4440/A1 U$$4347/A2 U$$4305/A1 U$$4347/B2 VGND VGND VPWR VPWR U$$4304/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4314 U$$4314/A U$$4334/B VGND VGND VPWR VPWR U$$4314/X sky130_fd_sc_hd__xor2_1
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4325 _587_/Q U$$4335/A2 _588_/Q U$$4333/B2 VGND VGND VPWR VPWR U$$4326/A sky130_fd_sc_hd__a22o_1
XFILLER_78_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4336 U$$4336/A _679_/Q VGND VGND VPWR VPWR U$$4336/X sky130_fd_sc_hd__xor2_1
XFILLER_133_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4347 U$$4484/A1 U$$4347/A2 U$$4486/A1 U$$4347/B2 VGND VGND VPWR VPWR U$$4348/A
+ sky130_fd_sc_hd__a22o_1
XU$$3602 U$$3602/A1 U$$3636/A2 U$$4426/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3603/A
+ sky130_fd_sc_hd__a22o_1
XU$$3613 U$$3613/A U$$3613/B VGND VGND VPWR VPWR U$$3613/X sky130_fd_sc_hd__xor2_1
XU$$4358 U$$4358/A U$$4382/B VGND VGND VPWR VPWR U$$4358/X sky130_fd_sc_hd__xor2_1
XFILLER_19_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3624 U$$3624/A1 U$$3662/A2 U$$4448/A1 U$$3662/B2 VGND VGND VPWR VPWR U$$3625/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4369 U$$4369/A1 U$$4369/A2 U$$4369/B1 U$$4369/B2 VGND VGND VPWR VPWR U$$4370/A
+ sky130_fd_sc_hd__a22o_1
XU$$3635 U$$3635/A U$$3637/B VGND VGND VPWR VPWR U$$3635/X sky130_fd_sc_hd__xor2_1
XU$$2901 U$$3175/A1 U$$2915/A2 U$$4410/A1 U$$2915/B2 VGND VGND VPWR VPWR U$$2902/A
+ sky130_fd_sc_hd__a22o_1
XU$$3646 U$$3646/A1 U$$3664/A2 U$$4470/A1 U$$3664/B2 VGND VGND VPWR VPWR U$$3647/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3657 U$$3657/A U$$3671/B VGND VGND VPWR VPWR U$$3657/X sky130_fd_sc_hd__xor2_1
XU$$2912 U$$2912/A U$$2966/B VGND VGND VPWR VPWR U$$2912/X sky130_fd_sc_hd__xor2_1
XU$$2923 U$$731/A1 U$$2929/A2 U$$596/A1 U$$2929/B2 VGND VGND VPWR VPWR U$$2924/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_108_2 dadda_fa_4_108_2/A dadda_fa_4_108_2/B dadda_fa_4_108_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/CIN dadda_fa_5_108_1/CIN sky130_fd_sc_hd__fa_1
XU$$3668 U$$3805/A1 U$$3566/X U$$3805/B1 U$$3567/X VGND VGND VPWR VPWR U$$3669/A sky130_fd_sc_hd__a22o_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2934 U$$2934/A U$$2972/B VGND VGND VPWR VPWR U$$2934/X sky130_fd_sc_hd__xor2_1
XFILLER_46_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3679 U$$3679/A U$$3698/A VGND VGND VPWR VPWR U$$3679/X sky130_fd_sc_hd__xor2_1
XU$$2945 U$$3493/A1 U$$2981/A2 U$$3495/A1 U$$2981/B2 VGND VGND VPWR VPWR U$$2946/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2956 U$$2956/A U$$2982/B VGND VGND VPWR VPWR U$$2956/X sky130_fd_sc_hd__xor2_1
XFILLER_61_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_250 _195_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2967 U$$4472/B1 U$$2881/X U$$4476/A1 U$$2882/X VGND VGND VPWR VPWR U$$2968/A sky130_fd_sc_hd__a22o_1
XANTENNA_261 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2978 U$$2978/A U$$2982/B VGND VGND VPWR VPWR U$$2978/X sky130_fd_sc_hd__xor2_1
XANTENNA_272 _199_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_508_ _516_/CLK _508_/D VGND VGND VPWR VPWR _508_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2989 U$$3124/B1 U$$2997/A2 U$$2991/A1 U$$2997/B2 VGND VGND VPWR VPWR U$$2990/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_283 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_294 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_439_ _439_/CLK _439_/D VGND VGND VPWR VPWR _439_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_clk _616_/CLK VGND VGND VPWR VPWR _486_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_81_2 dadda_fa_2_81_2/A dadda_fa_2_81_2/B dadda_fa_2_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/A dadda_fa_3_81_3/A sky130_fd_sc_hd__fa_1
XFILLER_115_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_74_1 dadda_fa_2_74_1/A dadda_fa_2_74_1/B dadda_fa_2_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_0/CIN dadda_fa_3_74_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_51_0 dadda_fa_5_51_0/A dadda_fa_5_51_0/B dadda_fa_5_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_52_0/A dadda_fa_6_51_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_67_0 dadda_fa_2_67_0/A dadda_fa_2_67_0/B dadda_fa_2_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_0/B dadda_fa_3_67_2/B sky130_fd_sc_hd__fa_1
XFILLER_68_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1057 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_31_clk _479_/CLK VGND VGND VPWR VPWR _475_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_96_2 dadda_fa_4_96_2/A dadda_fa_4_96_2/B dadda_fa_4_96_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/CIN dadda_fa_5_96_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_138_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_89_1 dadda_fa_4_89_1/A dadda_fa_4_89_1/B dadda_fa_4_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/B dadda_fa_5_89_1/B sky130_fd_sc_hd__fa_1
XFILLER_156_1112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_66_0 dadda_fa_7_66_0/A dadda_fa_7_66_0/B dadda_fa_7_66_0/CIN VGND VGND
+ VPWR VPWR _491_/D _362_/D sky130_fd_sc_hd__fa_1
XFILLER_69_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1025 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2208 U$$2345/A1 U$$2242/A2 U$$2895/A1 U$$2242/B2 VGND VGND VPWR VPWR U$$2209/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2219 U$$2219/A U$$2263/B VGND VGND VPWR VPWR U$$2219/X sky130_fd_sc_hd__xor2_1
XFILLER_170_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4385_1768 VGND VGND VPWR VPWR U$$4385_1768/HI U$$4385/A sky130_fd_sc_hd__conb_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1507 U$$1507/A VGND VGND VPWR VPWR U$$1507/Y sky130_fd_sc_hd__inv_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1518 U$$1518/A U$$1558/B VGND VGND VPWR VPWR U$$1518/X sky130_fd_sc_hd__xor2_1
XFILLER_76_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1529 U$$568/B1 U$$1557/A2 U$$435/A1 U$$1557/B2 VGND VGND VPWR VPWR U$$1530/A sky130_fd_sc_hd__a22o_1
XFILLER_103_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk _432_/CLK VGND VGND VPWR VPWR _428_/CLK sky130_fd_sc_hd__clkbuf_16
X_224_ _225_/CLK _224_/D VGND VGND VPWR VPWR _224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_91_1 dadda_fa_3_91_1/A dadda_fa_3_91_1/B dadda_fa_3_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_0/CIN dadda_fa_4_91_2/A sky130_fd_sc_hd__fa_1
XFILLER_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_84_0 dadda_fa_3_84_0/A dadda_fa_3_84_0/B dadda_fa_3_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_0/B dadda_fa_4_84_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_174_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_89_clk _628_/CLK VGND VGND VPWR VPWR _624_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater407 U$$689/X VGND VGND VPWR VPWR U$$795/A2 sky130_fd_sc_hd__buf_4
Xrepeater418 U$$4381/A2 VGND VGND VPWR VPWR U$$4369/A2 sky130_fd_sc_hd__buf_6
XU$$4100 U$$4100/A U$$4109/A VGND VGND VPWR VPWR U$$4100/X sky130_fd_sc_hd__xor2_1
XU$$4111 _676_/Q VGND VGND VPWR VPWR U$$4113/B sky130_fd_sc_hd__inv_1
Xrepeater429 U$$545/A2 VGND VGND VPWR VPWR U$$517/A2 sky130_fd_sc_hd__buf_4
XU$$4122 U$$4396/A1 U$$4140/A2 U$$4259/B1 U$$4140/B2 VGND VGND VPWR VPWR U$$4123/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4133 U$$4133/A U$$4215/B VGND VGND VPWR VPWR U$$4133/X sky130_fd_sc_hd__xor2_1
XU$$4144 U$$4418/A1 U$$4182/A2 U$$4418/B1 U$$4182/B2 VGND VGND VPWR VPWR U$$4145/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4155 U$$4155/A U$$4183/B VGND VGND VPWR VPWR U$$4155/X sky130_fd_sc_hd__xor2_1
XFILLER_66_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3410 U$$4506/A1 U$$3292/X U$$3412/A1 U$$3293/X VGND VGND VPWR VPWR U$$3411/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_113_0 U$$4223/X U$$4356/X U$$4489/X VGND VGND VPWR VPWR dadda_fa_5_114_0/A
+ dadda_fa_5_113_1/A sky130_fd_sc_hd__fa_1
XU$$3421 U$$3421/A U$$3423/B VGND VGND VPWR VPWR U$$3421/X sky130_fd_sc_hd__xor2_1
XU$$4166 U$$4440/A1 U$$4226/A2 U$$4305/A1 U$$4226/B2 VGND VGND VPWR VPWR U$$4167/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_46_5 dadda_fa_2_46_5/A dadda_fa_2_46_5/B dadda_fa_2_46_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_2/A dadda_fa_4_46_0/A sky130_fd_sc_hd__fa_1
XU$$3432 U$$3432/A U$$3478/B VGND VGND VPWR VPWR U$$3432/X sky130_fd_sc_hd__xor2_1
XU$$4177 U$$4177/A U$$4203/B VGND VGND VPWR VPWR U$$4177/X sky130_fd_sc_hd__xor2_1
XU$$4188 _587_/Q U$$4196/A2 _588_/Q U$$4196/B2 VGND VGND VPWR VPWR U$$4189/A sky130_fd_sc_hd__a22o_1
XU$$3443 U$$3578/B1 U$$3479/A2 U$$3445/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3444/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4199 U$$4199/A U$$4203/B VGND VGND VPWR VPWR U$$4199/X sky130_fd_sc_hd__xor2_1
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3454 U$$3454/A U$$3498/B VGND VGND VPWR VPWR U$$3454/X sky130_fd_sc_hd__xor2_1
XFILLER_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_39_4 input189/X dadda_fa_2_39_4/B dadda_fa_2_39_4/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_40_1/CIN dadda_fa_3_39_3/CIN sky130_fd_sc_hd__fa_1
XU$$2720 U$$2720/A U$$2730/B VGND VGND VPWR VPWR U$$2720/X sky130_fd_sc_hd__xor2_1
XU$$3465 U$$3602/A1 U$$3559/A2 U$$4426/A1 U$$3559/B2 VGND VGND VPWR VPWR U$$3466/A
+ sky130_fd_sc_hd__a22o_1
XU$$2731 U$$3005/A1 U$$2733/A2 _613_/Q U$$2733/B2 VGND VGND VPWR VPWR U$$2732/A sky130_fd_sc_hd__a22o_1
XU$$3476 U$$3476/A U$$3478/B VGND VGND VPWR VPWR U$$3476/X sky130_fd_sc_hd__xor2_1
XU$$3487 U$$3624/A1 U$$3519/A2 _580_/Q U$$3519/B2 VGND VGND VPWR VPWR U$$3488/A sky130_fd_sc_hd__a22o_1
XU$$2742 U$$2877/A VGND VGND VPWR VPWR U$$2742/Y sky130_fd_sc_hd__inv_1
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2753 U$$2753/A U$$2795/B VGND VGND VPWR VPWR U$$2753/X sky130_fd_sc_hd__xor2_1
XU$$3498 U$$3498/A U$$3498/B VGND VGND VPWR VPWR U$$3498/X sky130_fd_sc_hd__xor2_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2764 U$$981/B1 U$$2812/A2 U$$3312/B1 U$$2812/B2 VGND VGND VPWR VPWR U$$2765/A
+ sky130_fd_sc_hd__a22o_1
XU$$2775 U$$2775/A U$$2827/B VGND VGND VPWR VPWR U$$2775/X sky130_fd_sc_hd__xor2_1
XFILLER_178_215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2786 U$$731/A1 U$$2788/A2 U$$2786/B1 U$$2788/B2 VGND VGND VPWR VPWR U$$2787/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2797 U$$2797/A U$$2839/B VGND VGND VPWR VPWR U$$2797/X sky130_fd_sc_hd__xor2_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk _616_/CLK VGND VGND VPWR VPWR _470_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_99_0 dadda_fa_5_99_0/A dadda_fa_5_99_0/B dadda_fa_5_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_100_0/A dadda_fa_6_99_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$704 final_adder.U$$704/A final_adder.U$$704/B VGND VGND VPWR VPWR
+ _250_/D sky130_fd_sc_hd__xor2_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$715 final_adder.U$$715/A final_adder.U$$715/B VGND VGND VPWR VPWR
+ _261_/D sky130_fd_sc_hd__xor2_1
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$726 final_adder.U$$726/A final_adder.U$$726/B VGND VGND VPWR VPWR
+ _272_/D sky130_fd_sc_hd__xor2_4
Xrepeater930 _673_/Q VGND VGND VPWR VPWR U$$3973/A sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$737 final_adder.U$$737/A final_adder.U$$737/B VGND VGND VPWR VPWR
+ _283_/D sky130_fd_sc_hd__xor2_4
XFILLER_68_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater941 _671_/Q VGND VGND VPWR VPWR U$$3764/B sky130_fd_sc_hd__buf_6
XFILLER_25_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$748 final_adder.U$$748/A final_adder.U$$748/B VGND VGND VPWR VPWR
+ _294_/D sky130_fd_sc_hd__xor2_4
Xrepeater952 _669_/Q VGND VGND VPWR VPWR U$$3675/B sky130_fd_sc_hd__buf_6
XFILLER_112_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater963 U$$3538/B VGND VGND VPWR VPWR U$$3520/B sky130_fd_sc_hd__buf_8
XU$$609 U$$609/A U$$613/B VGND VGND VPWR VPWR U$$609/X sky130_fd_sc_hd__xor2_1
XFILLER_72_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater974 _665_/Q VGND VGND VPWR VPWR U$$3425/A sky130_fd_sc_hd__buf_6
Xrepeater985 U$$3077/B VGND VGND VPWR VPWR U$$3049/B sky130_fd_sc_hd__buf_8
Xrepeater996 U$$2982/B VGND VGND VPWR VPWR U$$2966/B sky130_fd_sc_hd__buf_12
XFILLER_186_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_90_0_1859 VGND VGND VPWR VPWR dadda_fa_1_90_0/A dadda_fa_1_90_0_1859/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1509 U$$467/A1 VGND VGND VPWR VPWR U$$878/A1 sky130_fd_sc_hd__buf_4
XFILLER_158_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_108_1 U$$3681/X U$$3814/X U$$3947/X VGND VGND VPWR VPWR dadda_fa_4_109_0/CIN
+ dadda_fa_4_108_2/A sky130_fd_sc_hd__fa_1
XFILLER_109_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput290 _182_/Q VGND VGND VPWR VPWR o[14] sky130_fd_sc_hd__buf_2
XFILLER_43_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_49_3 dadda_fa_3_49_3/A dadda_fa_3_49_3/B dadda_fa_3_49_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_1/B dadda_fa_4_49_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2005 U$$2005/A U$$2043/B VGND VGND VPWR VPWR U$$2005/X sky130_fd_sc_hd__xor2_1
XFILLER_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2016 U$$781/B1 U$$2028/A2 U$$3386/B1 U$$2028/B2 VGND VGND VPWR VPWR U$$2017/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2027 U$$2027/A U$$2054/A VGND VGND VPWR VPWR U$$2027/X sky130_fd_sc_hd__xor2_1
XU$$2038 U$$940/B1 U$$2038/A2 U$$944/A1 U$$2038/B2 VGND VGND VPWR VPWR U$$2039/A sky130_fd_sc_hd__a22o_1
XU$$1304 U$$1304/A U$$1310/B VGND VGND VPWR VPWR U$$1304/X sky130_fd_sc_hd__xor2_1
XU$$2049 U$$2049/A U$$2054/A VGND VGND VPWR VPWR U$$2049/X sky130_fd_sc_hd__xor2_1
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1315 U$$3096/A1 U$$1355/A2 U$$3096/B1 U$$1355/B2 VGND VGND VPWR VPWR U$$1316/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1326 U$$1326/A U$$1332/B VGND VGND VPWR VPWR U$$1326/X sky130_fd_sc_hd__xor2_1
XFILLER_43_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1337 U$$926/A1 U$$1237/X U$$928/A1 U$$1238/X VGND VGND VPWR VPWR U$$1338/A sky130_fd_sc_hd__a22o_1
XFILLER_16_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1348 U$$1348/A U$$1356/B VGND VGND VPWR VPWR U$$1348/X sky130_fd_sc_hd__xor2_1
XFILLER_200_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1359 U$$948/A1 U$$1367/A2 _612_/Q U$$1367/B2 VGND VGND VPWR VPWR U$$1360/A sky130_fd_sc_hd__a22o_1
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_207_ _207_/CLK _207_/D VGND VGND VPWR VPWR _207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_808 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_616 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_2_clk _442_/CLK VGND VGND VPWR VPWR _443_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_51_3 dadda_fa_2_51_3/A dadda_fa_2_51_3/B dadda_fa_2_51_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/B dadda_fa_3_51_3/B sky130_fd_sc_hd__fa_1
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_44_2 U$$3065/B input195/X dadda_fa_2_44_2/CIN VGND VGND VPWR VPWR dadda_fa_3_45_1/A
+ dadda_fa_3_44_3/A sky130_fd_sc_hd__fa_1
XFILLER_65_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$11 _435_/Q _307_/Q VGND VGND VPWR VPWR final_adder.U$$139/B1 final_adder.U$$633/A
+ sky130_fd_sc_hd__ha_2
XU$$3240 U$$3240/A U$$3286/B VGND VGND VPWR VPWR U$$3240/X sky130_fd_sc_hd__xor2_1
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_21_1 dadda_fa_5_21_1/A dadda_fa_5_21_1/B dadda_fa_5_21_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_22_0/B dadda_fa_7_21_0/A sky130_fd_sc_hd__fa_1
XU$$3251 U$$3386/B1 U$$3263/A2 U$$3388/B1 U$$3263/B2 VGND VGND VPWR VPWR U$$3252/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$22 _446_/Q _318_/Q VGND VGND VPWR VPWR final_adder.U$$517/B1 final_adder.U$$644/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$33 _457_/Q _329_/Q VGND VGND VPWR VPWR final_adder.U$$161/B1 final_adder.U$$655/A
+ sky130_fd_sc_hd__ha_1
XU$$3262 U$$3262/A U$$3272/B VGND VGND VPWR VPWR U$$3262/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_37_1 U$$1145/X U$$1278/X U$$1411/X VGND VGND VPWR VPWR dadda_fa_3_38_0/CIN
+ dadda_fa_3_37_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$44 _468_/Q _340_/Q VGND VGND VPWR VPWR final_adder.U$$539/B1 final_adder.U$$666/A
+ sky130_fd_sc_hd__ha_2
XU$$3273 U$$3273/A1 U$$3273/A2 U$$3412/A1 U$$3273/B2 VGND VGND VPWR VPWR U$$3274/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$55 _479_/Q _351_/Q VGND VGND VPWR VPWR final_adder.U$$183/B1 final_adder.U$$677/A
+ sky130_fd_sc_hd__ha_1
XFILLER_53_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_14_0 dadda_fa_5_14_0/A dadda_fa_5_14_0/B dadda_fa_5_14_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_15_0/A dadda_fa_6_14_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3284 U$$3284/A U$$3288/A VGND VGND VPWR VPWR U$$3284/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$66 _490_/Q _362_/Q VGND VGND VPWR VPWR final_adder.U$$561/B1 final_adder.U$$688/A
+ sky130_fd_sc_hd__ha_2
XU$$2550 U$$906/A1 U$$2550/A2 U$$908/A1 U$$2550/B2 VGND VGND VPWR VPWR U$$2551/A sky130_fd_sc_hd__a22o_1
XFILLER_62_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3295 U$$3295/A U$$3343/B VGND VGND VPWR VPWR U$$3295/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$77 _501_/Q _373_/Q VGND VGND VPWR VPWR final_adder.U$$205/B1 final_adder.U$$699/A
+ sky130_fd_sc_hd__ha_1
XU$$2561 U$$2561/A U$$2567/B VGND VGND VPWR VPWR U$$2561/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2572 U$$4353/A1 U$$2580/A2 U$$4490/B1 U$$2580/B2 VGND VGND VPWR VPWR U$$2573/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$88 _512_/Q _384_/Q VGND VGND VPWR VPWR final_adder.U$$583/B1 final_adder.U$$710/A
+ sky130_fd_sc_hd__ha_2
XFILLER_206_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$99 _523_/Q _395_/Q VGND VGND VPWR VPWR final_adder.U$$227/B1 final_adder.U$$721/A
+ sky130_fd_sc_hd__ha_1
XFILLER_179_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2583 U$$2583/A U$$2583/B VGND VGND VPWR VPWR U$$2583/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2594 _612_/Q U$$2600/A2 _613_/Q U$$2600/B2 VGND VGND VPWR VPWR U$$2595/A sky130_fd_sc_hd__a22o_1
XFILLER_21_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1860 U$$1860/A U$$1870/B VGND VGND VPWR VPWR U$$1860/X sky130_fd_sc_hd__xor2_1
XFILLER_34_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1871 U$$4474/A1 U$$1907/A2 U$$3380/A1 U$$1907/B2 VGND VGND VPWR VPWR U$$1872/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1882 U$$1882/A U$$1884/B VGND VGND VPWR VPWR U$$1882/X sky130_fd_sc_hd__xor2_1
XU$$1893 U$$384/B1 U$$1897/A2 U$$251/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1894/A sky130_fd_sc_hd__a22o_1
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_1_40_3 U$$1284/X U$$1417/X VGND VGND VPWR VPWR dadda_fa_2_41_4/CIN dadda_fa_3_40_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_118_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_59_2 dadda_fa_4_59_2/A dadda_fa_4_59_2/B dadda_fa_4_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/CIN dadda_fa_5_59_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$501 final_adder.U$$628/A final_adder.U$$628/B final_adder.U$$6/COUT
+ VGND VGND VPWR VPWR final_adder.U$$629/B sky130_fd_sc_hd__a21o_1
XTAP_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$523 final_adder.U$$650/A final_adder.U$$650/B final_adder.U$$523/B1
+ VGND VGND VPWR VPWR final_adder.U$$651/B sky130_fd_sc_hd__a21o_1
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_4_10_1 U$$426/X U$$559/X VGND VGND VPWR VPWR dadda_fa_5_11_1/A dadda_ha_4_10_1/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_85_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$545 final_adder.U$$672/A final_adder.U$$672/B final_adder.U$$545/B1
+ VGND VGND VPWR VPWR final_adder.U$$673/B sky130_fd_sc_hd__a21o_1
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_29_0 dadda_fa_7_29_0/A dadda_fa_7_29_0/B dadda_fa_7_29_0/CIN VGND VGND
+ VPWR VPWR _454_/D _325_/D sky130_fd_sc_hd__fa_1
Xrepeater760 U$$2943/B2 VGND VGND VPWR VPWR U$$2915/B2 sky130_fd_sc_hd__buf_4
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$567 final_adder.U$$694/A final_adder.U$$694/B final_adder.U$$567/B1
+ VGND VGND VPWR VPWR final_adder.U$$695/B sky130_fd_sc_hd__a21o_1
XFILLER_29_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$406 U$$406/A1 U$$278/X U$$406/B1 U$$279/X VGND VGND VPWR VPWR U$$407/A sky130_fd_sc_hd__a22o_1
Xrepeater771 U$$392/B2 VGND VGND VPWR VPWR U$$350/B2 sky130_fd_sc_hd__buf_4
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$417 U$$417/A1 U$$447/A2 U$$8/A1 U$$447/B2 VGND VGND VPWR VPWR U$$418/A sky130_fd_sc_hd__a22o_1
Xrepeater782 U$$2745/X VGND VGND VPWR VPWR U$$2874/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$589 final_adder.U$$716/A final_adder.U$$716/B final_adder.U$$589/B1
+ VGND VGND VPWR VPWR final_adder.U$$717/B sky130_fd_sc_hd__a21o_1
XFILLER_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$428 U$$428/A U$$456/B VGND VGND VPWR VPWR U$$428/X sky130_fd_sc_hd__xor2_1
Xrepeater793 U$$2524/B2 VGND VGND VPWR VPWR U$$2516/B2 sky130_fd_sc_hd__buf_4
XU$$439 U$$28/A1 U$$457/A2 U$$30/A1 U$$457/B2 VGND VGND VPWR VPWR U$$440/A sky130_fd_sc_hd__a22o_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1306 U$$791/A1 VGND VGND VPWR VPWR U$$515/B1 sky130_fd_sc_hd__buf_6
XFILLER_10_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1317 _600_/Q VGND VGND VPWR VPWR U$$3253/B1 sky130_fd_sc_hd__buf_4
Xrepeater1328 U$$4486/A1 VGND VGND VPWR VPWR U$$2705/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_107_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1339 U$$3521/B1 VGND VGND VPWR VPWR U$$98/A1 sky130_fd_sc_hd__buf_6
XFILLER_153_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_61_2 dadda_fa_3_61_2/A dadda_fa_3_61_2/B dadda_fa_3_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_1/A dadda_fa_4_61_2/B sky130_fd_sc_hd__fa_1
XFILLER_95_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_54_1 dadda_fa_3_54_1/A dadda_fa_3_54_1/B dadda_fa_3_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_0/CIN dadda_fa_4_54_2/A sky130_fd_sc_hd__fa_1
XFILLER_0_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_31_0 dadda_fa_6_31_0/A dadda_fa_6_31_0/B dadda_fa_6_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_32_0/B dadda_fa_7_31_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_47_0 dadda_fa_3_47_0/A dadda_fa_3_47_0/B dadda_fa_3_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_0/B dadda_fa_4_47_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$940 U$$940/A1 U$$948/A2 U$$940/B1 U$$948/B2 VGND VGND VPWR VPWR U$$941/A sky130_fd_sc_hd__a22o_1
XU$$951 U$$951/A U$$951/B VGND VGND VPWR VPWR U$$951/X sky130_fd_sc_hd__xor2_1
XU$$962 _631_/Q U$$962/B VGND VGND VPWR VPWR U$$962/X sky130_fd_sc_hd__and2_1
XU$$1101 U$$1099/B _631_/Q _632_/Q U$$1096/Y VGND VGND VPWR VPWR U$$1101/X sky130_fd_sc_hd__a22o_1
XFILLER_90_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1112 U$$16/A1 U$$1146/A2 U$$18/A1 U$$1146/B2 VGND VGND VPWR VPWR U$$1113/A sky130_fd_sc_hd__a22o_1
XFILLER_16_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$973 U$$973/A1 U$$995/A2 U$$973/B1 U$$995/B2 VGND VGND VPWR VPWR U$$974/A sky130_fd_sc_hd__a22o_1
XU$$1123 U$$1123/A U$$1151/B VGND VGND VPWR VPWR U$$1123/X sky130_fd_sc_hd__xor2_1
XFILLER_90_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$984 U$$984/A U$$998/B VGND VGND VPWR VPWR U$$984/X sky130_fd_sc_hd__xor2_1
XFILLER_188_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1134 U$$449/A1 U$$1146/A2 U$$449/B1 U$$1146/B2 VGND VGND VPWR VPWR U$$1135/A sky130_fd_sc_hd__a22o_1
XU$$995 U$$36/A1 U$$995/A2 U$$38/A1 U$$995/B2 VGND VGND VPWR VPWR U$$996/A sky130_fd_sc_hd__a22o_1
XFILLER_31_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1145 U$$1145/A U$$1147/B VGND VGND VPWR VPWR U$$1145/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1156 U$$60/A1 U$$1190/A2 U$$62/A1 U$$1190/B2 VGND VGND VPWR VPWR U$$1157/A sky130_fd_sc_hd__a22o_1
XU$$1167 U$$1167/A U$$1177/B VGND VGND VPWR VPWR U$$1167/X sky130_fd_sc_hd__xor2_1
XU$$1178 U$$80/B1 U$$1224/A2 U$$906/A1 U$$1224/B2 VGND VGND VPWR VPWR U$$1179/A sky130_fd_sc_hd__a22o_1
XFILLER_43_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1189 U$$1189/A U$$1209/B VGND VGND VPWR VPWR U$$1189/X sky130_fd_sc_hd__xor2_1
XFILLER_203_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_104_0 dadda_fa_7_104_0/A dadda_fa_7_104_0/B dadda_fa_7_104_0/CIN VGND
+ VGND VPWR VPWR _529_/D _400_/D sky130_fd_sc_hd__fa_1
XFILLER_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_99_3 U$$3663/X U$$3796/X U$$3929/X VGND VGND VPWR VPWR dadda_fa_3_100_2/A
+ dadda_fa_3_99_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_5_69_1 dadda_fa_5_69_1/A dadda_fa_5_69_1/B dadda_fa_5_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_70_0/B dadda_fa_7_69_0/A sky130_fd_sc_hd__fa_2
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3070 U$$4301/B1 U$$3148/A2 U$$4305/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3071/A
+ sky130_fd_sc_hd__a22o_1
XU$$3081 U$$3081/A U$$3083/B VGND VGND VPWR VPWR U$$3081/X sky130_fd_sc_hd__xor2_1
XU$$3092 U$$4051/A1 U$$3120/A2 U$$4053/A1 U$$3120/B2 VGND VGND VPWR VPWR U$$3093/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2380 U$$2380/A U$$2436/B VGND VGND VPWR VPWR U$$2380/X sky130_fd_sc_hd__xor2_1
XFILLER_210_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2391 U$$334/B1 U$$2395/A2 U$$64/A1 U$$2395/B2 VGND VGND VPWR VPWR U$$2392/A sky130_fd_sc_hd__a22o_1
XFILLER_22_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1690 U$$731/A1 U$$1740/A2 U$$733/A1 U$$1740/B2 VGND VGND VPWR VPWR U$$1691/A sky130_fd_sc_hd__a22o_1
XFILLER_210_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_71_1 dadda_fa_4_71_1/A dadda_fa_4_71_1/B dadda_fa_4_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/B dadda_fa_5_71_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_87_1 U$$2043/X U$$2176/X U$$2309/X VGND VGND VPWR VPWR dadda_fa_2_88_3/B
+ dadda_fa_2_87_5/A sky130_fd_sc_hd__fa_1
XFILLER_89_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_64_0 dadda_fa_4_64_0/A dadda_fa_4_64_0/B dadda_fa_4_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/A dadda_fa_5_64_1/A sky130_fd_sc_hd__fa_1
XTAP_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_610_ _613_/CLK _610_/D VGND VGND VPWR VPWR _610_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$331 final_adder.U$$330/A final_adder.U$$277/X final_adder.U$$279/X
+ VGND VGND VPWR VPWR final_adder.U$$331/X sky130_fd_sc_hd__a21o_1
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$342 final_adder.U$$342/A final_adder.U$$342/B VGND VGND VPWR VPWR
+ final_adder.U$$362/A sky130_fd_sc_hd__and2_1
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$353 final_adder.U$$322/X final_adder.U$$630/B final_adder.U$$323/X
+ VGND VGND VPWR VPWR final_adder.U$$638/B sky130_fd_sc_hd__a21o_4
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$364 final_adder.U$$364/A final_adder.U$$364/B VGND VGND VPWR VPWR
+ final_adder.U$$364/X sky130_fd_sc_hd__and2_1
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_934 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$203 U$$614/A1 U$$217/A2 U$$614/B1 U$$217/B2 VGND VGND VPWR VPWR U$$204/A sky130_fd_sc_hd__a22o_1
XFILLER_176_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$214 U$$214/A U$$216/B VGND VGND VPWR VPWR U$$214/X sky130_fd_sc_hd__xor2_1
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_541_ _541_/CLK _541_/D VGND VGND VPWR VPWR _541_/Q sky130_fd_sc_hd__dfxtp_1
XU$$225 U$$88/A1 U$$263/A2 U$$90/A1 U$$263/B2 VGND VGND VPWR VPWR U$$226/A sky130_fd_sc_hd__a22o_1
Xrepeater590 U$$1785/X VGND VGND VPWR VPWR U$$1907/A2 sky130_fd_sc_hd__buf_8
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$397 final_adder.U$$360/B final_adder.U$$686/B final_adder.U$$337/X
+ VGND VGND VPWR VPWR final_adder.U$$694/B sky130_fd_sc_hd__a21o_2
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$236 U$$236/A U$$250/B VGND VGND VPWR VPWR U$$236/X sky130_fd_sc_hd__xor2_1
XU$$247 U$$382/B1 U$$249/A2 U$$384/B1 U$$249/B2 VGND VGND VPWR VPWR U$$248/A sky130_fd_sc_hd__a22o_1
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$258 U$$258/A U$$264/B VGND VGND VPWR VPWR U$$258/X sky130_fd_sc_hd__xor2_1
XU$$269 U$$406/A1 U$$141/X U$$406/B1 U$$142/X VGND VGND VPWR VPWR U$$270/A sky130_fd_sc_hd__a22o_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_472_ _476_/CLK _472_/D VGND VGND VPWR VPWR _472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_499 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$8 U$$8/A1 U$$8/A2 U$$8/B1 U$$8/B2 VGND VGND VPWR VPWR U$$9/A sky130_fd_sc_hd__a22o_1
Xrepeater1103 U$$1296/B VGND VGND VPWR VPWR U$$1280/B sky130_fd_sc_hd__buf_6
XFILLER_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1114 U$$1203/B VGND VGND VPWR VPWR U$$1191/B sky130_fd_sc_hd__buf_6
Xdadda_ha_0_76_1 U$$1223/X U$$1356/X VGND VGND VPWR VPWR dadda_fa_1_77_8/CIN dadda_fa_2_76_0/A
+ sky130_fd_sc_hd__ha_1
Xrepeater1125 U$$1078/B VGND VGND VPWR VPWR U$$998/B sky130_fd_sc_hd__buf_8
Xdadda_fa_6_79_0 dadda_fa_6_79_0/A dadda_fa_6_79_0/B dadda_fa_6_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_80_0/B dadda_fa_7_79_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1136 U$$935/B VGND VGND VPWR VPWR U$$951/B sky130_fd_sc_hd__buf_12
Xrepeater1147 U$$659/B VGND VGND VPWR VPWR U$$613/B sky130_fd_sc_hd__clkbuf_8
XFILLER_153_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1158 U$$500/B VGND VGND VPWR VPWR U$$484/B sky130_fd_sc_hd__buf_6
XFILLER_153_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1169 U$$410/A VGND VGND VPWR VPWR U$$383/B sky130_fd_sc_hd__buf_6
XFILLER_141_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_411 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$770 U$$770/A U$$816/B VGND VGND VPWR VPWR U$$770/X sky130_fd_sc_hd__xor2_1
XFILLER_1_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$781 U$$916/B1 U$$783/A2 U$$781/B1 U$$783/B2 VGND VGND VPWR VPWR U$$782/A sky130_fd_sc_hd__a22o_1
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$792 U$$792/A U$$810/B VGND VGND VPWR VPWR U$$792/X sky130_fd_sc_hd__xor2_1
XFILLER_44_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_81_0 dadda_fa_5_81_0/A dadda_fa_5_81_0/B dadda_fa_5_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_82_0/A dadda_fa_6_81_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_97_0 U$$2328/Y U$$2462/X U$$2595/X VGND VGND VPWR VPWR dadda_fa_3_98_0/B
+ dadda_fa_3_97_2/B sky130_fd_sc_hd__fa_1
XFILLER_172_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1670 _557_/Q VGND VGND VPWR VPWR U$$3578/B1 sky130_fd_sc_hd__buf_6
Xrepeater1681 U$$2754/A1 VGND VGND VPWR VPWR U$$973/A1 sky130_fd_sc_hd__buf_6
XFILLER_67_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1692 U$$3437/A1 VGND VGND VPWR VPWR U$$2478/A1 sky130_fd_sc_hd__buf_6
XFILLER_141_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_73_7 dadda_fa_1_73_7/A dadda_fa_1_73_7/B dadda_fa_1_73_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_74_2/CIN dadda_fa_2_73_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_66_6 dadda_fa_1_66_6/A dadda_fa_1_66_6/B dadda_fa_1_66_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_2/B dadda_fa_2_66_5/B sky130_fd_sc_hd__fa_1
XFILLER_73_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_59_5 U$$3583/X U$$3716/X U$$3849/X VGND VGND VPWR VPWR dadda_fa_2_60_2/A
+ dadda_fa_2_59_5/A sky130_fd_sc_hd__fa_1
XFILLER_27_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1041 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_455 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_96_0 dadda_fa_7_96_0/A dadda_fa_7_96_0/B dadda_fa_7_96_0/CIN VGND VGND
+ VPWR VPWR _521_/D _392_/D sky130_fd_sc_hd__fa_1
XFILLER_183_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1222 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_23 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4507 U$$4507/A U$$4507/B VGND VGND VPWR VPWR U$$4507/X sky130_fd_sc_hd__xor2_1
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_111_0 dadda_fa_6_111_0/A dadda_fa_6_111_0/B dadda_fa_6_111_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_112_0/B dadda_fa_7_111_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1040 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3806 U$$3806/A _671_/Q VGND VGND VPWR VPWR U$$3806/X sky130_fd_sc_hd__xor2_1
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3817 U$$3952/B1 U$$3703/X U$$4504/A1 U$$3704/X VGND VGND VPWR VPWR U$$3818/A sky130_fd_sc_hd__a22o_1
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3828 U$$3828/A U$$3832/B VGND VGND VPWR VPWR U$$3828/X sky130_fd_sc_hd__xor2_1
XFILLER_18_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$150 final_adder.U$$645/A final_adder.U$$644/A VGND VGND VPWR VPWR
+ final_adder.U$$266/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$161 final_adder.U$$655/A final_adder.U$$527/B1 final_adder.U$$161/B1
+ VGND VGND VPWR VPWR final_adder.U$$161/X sky130_fd_sc_hd__a21o_1
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$172 final_adder.U$$667/A final_adder.U$$666/A VGND VGND VPWR VPWR
+ final_adder.U$$278/B sky130_fd_sc_hd__and2_1
XU$$3839 _673_/Q U$$3839/B VGND VGND VPWR VPWR U$$3839/X sky130_fd_sc_hd__and2_1
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_3 dadda_fa_3_31_3/A dadda_fa_3_31_3/B dadda_fa_3_31_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_1/B dadda_fa_4_31_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$183 final_adder.U$$677/A final_adder.U$$549/B1 final_adder.U$$183/B1
+ VGND VGND VPWR VPWR final_adder.U$$183/X sky130_fd_sc_hd__a21o_1
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$194 final_adder.U$$689/A final_adder.U$$688/A VGND VGND VPWR VPWR
+ final_adder.U$$288/A sky130_fd_sc_hd__and2_1
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_524_ _526_/CLK _524_/D VGND VGND VPWR VPWR _524_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_24_2 U$$1518/X U$$1651/X U$$1723/B VGND VGND VPWR VPWR dadda_fa_4_25_1/A
+ dadda_fa_4_24_2/B sky130_fd_sc_hd__fa_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_455_ _455_/CLK _455_/D VGND VGND VPWR VPWR _455_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_386_ _558_/CLK _386_/D VGND VGND VPWR VPWR _386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_76_5 dadda_fa_2_76_5/A dadda_fa_2_76_5/B dadda_fa_2_76_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_2/A dadda_fa_4_76_0/A sky130_fd_sc_hd__fa_1
XFILLER_141_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_69_4 dadda_fa_2_69_4/A dadda_fa_2_69_4/B dadda_fa_2_69_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/CIN dadda_fa_3_69_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_110_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput190 c[3] VGND VGND VPWR VPWR input190/X sky130_fd_sc_hd__clkbuf_4
XFILLER_3_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_444 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_106_1 dadda_fa_5_106_1/A dadda_fa_5_106_1/B dadda_fa_5_106_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_107_0/B dadda_fa_7_106_0/A sky130_fd_sc_hd__fa_2
XFILLER_145_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1010 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_71_4 U$$3740/X U$$3873/X U$$4006/X VGND VGND VPWR VPWR dadda_fa_2_72_1/CIN
+ dadda_fa_2_71_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_141_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_64_3 U$$3726/X U$$3859/X U$$3992/X VGND VGND VPWR VPWR dadda_fa_2_65_1/B
+ dadda_fa_2_64_4/B sky130_fd_sc_hd__fa_1
XFILLER_100_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_41_2 dadda_fa_4_41_2/A dadda_fa_4_41_2/B dadda_fa_4_41_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/CIN dadda_fa_5_41_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_57_2 U$$1983/X U$$2116/X U$$2249/X VGND VGND VPWR VPWR dadda_fa_2_58_1/A
+ dadda_fa_2_57_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_34_1 dadda_fa_4_34_1/A dadda_fa_4_34_1/B dadda_fa_4_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/B dadda_fa_5_34_1/B sky130_fd_sc_hd__fa_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_455 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_11_0 dadda_fa_7_11_0/A dadda_fa_7_11_0/B dadda_fa_7_11_0/CIN VGND VGND
+ VPWR VPWR _436_/D _307_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_27_0 dadda_fa_4_27_0/A dadda_fa_4_27_0/B dadda_fa_4_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/A dadda_fa_5_27_1/A sky130_fd_sc_hd__fa_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_240_ _372_/CLK _240_/D VGND VGND VPWR VPWR _240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_171_ _179_/CLK _171_/D VGND VGND VPWR VPWR _171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_0_60_4 U$$1723/X U$$1856/X VGND VGND VPWR VPWR dadda_fa_1_61_7/B dadda_fa_2_60_0/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_3_79_3 dadda_fa_3_79_3/A dadda_fa_3_79_3/B dadda_fa_3_79_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_1/B dadda_fa_4_79_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4304 U$$4304/A U$$4348/B VGND VGND VPWR VPWR U$$4304/X sky130_fd_sc_hd__xor2_1
XU$$4315 U$$4450/B1 U$$4327/A2 _583_/Q U$$4319/B2 VGND VGND VPWR VPWR U$$4316/A sky130_fd_sc_hd__a22o_1
XU$$4326 U$$4326/A U$$4334/B VGND VGND VPWR VPWR U$$4326/X sky130_fd_sc_hd__xor2_1
XU$$4337 U$$4472/B1 U$$4251/X U$$4337/B1 U$$4345/B2 VGND VGND VPWR VPWR U$$4338/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4348 U$$4348/A U$$4348/B VGND VGND VPWR VPWR U$$4348/X sky130_fd_sc_hd__xor2_1
XU$$3603 U$$3603/A U$$3637/B VGND VGND VPWR VPWR U$$3603/X sky130_fd_sc_hd__xor2_1
XFILLER_93_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3614 U$$3751/A1 U$$3662/A2 U$$3753/A1 U$$3662/B2 VGND VGND VPWR VPWR U$$3615/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4359 U$$934/A1 U$$4369/A2 U$$4498/A1 U$$4369/B2 VGND VGND VPWR VPWR U$$4360/A
+ sky130_fd_sc_hd__a22o_1
XU$$3625 U$$3625/A U$$3627/B VGND VGND VPWR VPWR U$$3625/X sky130_fd_sc_hd__xor2_1
XFILLER_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3636 U$$3771/B1 U$$3636/A2 U$$3638/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3637/A
+ sky130_fd_sc_hd__a22o_1
XU$$2902 U$$2902/A U$$2916/B VGND VGND VPWR VPWR U$$2902/X sky130_fd_sc_hd__xor2_1
XU$$3647 U$$3647/A U$$3663/B VGND VGND VPWR VPWR U$$3647/X sky130_fd_sc_hd__xor2_1
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2913 U$$719/B1 U$$2915/A2 U$$3187/B1 U$$2915/B2 VGND VGND VPWR VPWR U$$2914/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3658 U$$3658/A1 U$$3664/A2 _597_/Q U$$3664/B2 VGND VGND VPWR VPWR U$$3659/A sky130_fd_sc_hd__a22o_1
XFILLER_93_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2924 U$$2924/A U$$2928/B VGND VGND VPWR VPWR U$$2924/X sky130_fd_sc_hd__xor2_1
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3669 U$$3669/A U$$3671/B VGND VGND VPWR VPWR U$$3669/X sky130_fd_sc_hd__xor2_1
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2935 U$$4305/A1 U$$2973/A2 U$$4168/B1 U$$2973/B2 VGND VGND VPWR VPWR U$$2936/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2946 U$$2946/A U$$2966/B VGND VGND VPWR VPWR U$$2946/X sky130_fd_sc_hd__xor2_1
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_240 _192_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2957 U$$2957/A1 U$$2959/A2 U$$3916/B1 U$$2959/B2 VGND VGND VPWR VPWR U$$2958/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2968 U$$2968/A U$$3008/B VGND VGND VPWR VPWR U$$2968/X sky130_fd_sc_hd__xor2_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 _195_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_507_ _507_/CLK _507_/D VGND VGND VPWR VPWR _507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_262 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2979 U$$3799/B1 U$$3005/A2 U$$3529/A1 U$$3005/B2 VGND VGND VPWR VPWR U$$2980/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_273 _212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_284 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_295 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_438_ _439_/CLK _438_/D VGND VGND VPWR VPWR _438_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_369_ _369_/CLK _369_/D VGND VGND VPWR VPWR _369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_338 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$691_1843 VGND VGND VPWR VPWR U$$691_1843/HI U$$691/A1 sky130_fd_sc_hd__conb_1
XFILLER_154_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_81_3 dadda_fa_2_81_3/A dadda_fa_2_81_3/B dadda_fa_2_81_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/B dadda_fa_3_81_3/B sky130_fd_sc_hd__fa_1
XFILLER_103_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_74_2 dadda_fa_2_74_2/A dadda_fa_2_74_2/B dadda_fa_2_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/A dadda_fa_3_74_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_51_1 dadda_fa_5_51_1/A dadda_fa_5_51_1/B dadda_fa_5_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_52_0/B dadda_fa_7_51_0/A sky130_fd_sc_hd__fa_1
XFILLER_190_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_67_1 dadda_fa_2_67_1/A dadda_fa_2_67_1/B dadda_fa_2_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_0/CIN dadda_fa_3_67_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_44_0 dadda_fa_5_44_0/A dadda_fa_5_44_0/B dadda_fa_5_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_45_0/A dadda_fa_6_44_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_970 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_89_2 dadda_fa_4_89_2/A dadda_fa_4_89_2/B dadda_fa_4_89_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/CIN dadda_fa_5_89_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_59_0 dadda_fa_7_59_0/A dadda_fa_7_59_0/B dadda_fa_7_59_0/CIN VGND VGND
+ VPWR VPWR _484_/D _355_/D sky130_fd_sc_hd__fa_1
XFILLER_161_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_62_0 U$$2392/X U$$2525/X U$$2658/X VGND VGND VPWR VPWR dadda_fa_2_63_0/B
+ dadda_fa_2_62_3/B sky130_fd_sc_hd__fa_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_336 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2209 U$$2209/A U$$2241/B VGND VGND VPWR VPWR U$$2209/X sky130_fd_sc_hd__xor2_1
XFILLER_41_1084 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1508 _638_/Q VGND VGND VPWR VPWR U$$1510/B sky130_fd_sc_hd__inv_1
XFILLER_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1519 U$$2613/B1 U$$1557/A2 U$$2754/A1 U$$1557/B2 VGND VGND VPWR VPWR U$$1520/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_223_ _225_/CLK _223_/D VGND VGND VPWR VPWR _223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_91_2 dadda_fa_3_91_2/A dadda_fa_3_91_2/B dadda_fa_3_91_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_1/A dadda_fa_4_91_2/B sky130_fd_sc_hd__fa_1
XFILLER_48_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_84_1 dadda_fa_3_84_1/A dadda_fa_3_84_1/B dadda_fa_3_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_0/CIN dadda_fa_4_84_2/A sky130_fd_sc_hd__fa_1
XFILLER_128_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_61_0 dadda_fa_6_61_0/A dadda_fa_6_61_0/B dadda_fa_6_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_62_0/B dadda_fa_7_61_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_77_0 dadda_fa_3_77_0/A dadda_fa_3_77_0/B dadda_fa_3_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_0/B dadda_fa_4_77_1/CIN sky130_fd_sc_hd__fa_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater408 U$$689/X VGND VGND VPWR VPWR U$$809/A2 sky130_fd_sc_hd__buf_6
XU$$4101 U$$4512/A1 U$$4107/A2 U$$4514/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4102/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater419 U$$4251/X VGND VGND VPWR VPWR U$$4381/A2 sky130_fd_sc_hd__buf_4
XFILLER_144_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4112 _677_/Q VGND VGND VPWR VPWR U$$4112/Y sky130_fd_sc_hd__inv_1
XU$$4123 U$$4123/A U$$4141/B VGND VGND VPWR VPWR U$$4123/X sky130_fd_sc_hd__xor2_1
XU$$4134 U$$4408/A1 U$$4174/A2 U$$4273/A1 U$$4174/B2 VGND VGND VPWR VPWR U$$4135/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4145 U$$4145/A U$$4183/B VGND VGND VPWR VPWR U$$4145/X sky130_fd_sc_hd__xor2_1
XU$$3400 _604_/Q U$$3402/A2 U$$3539/A1 U$$3402/B2 VGND VGND VPWR VPWR U$$3401/A sky130_fd_sc_hd__a22o_1
XU$$4156 _571_/Q U$$4182/A2 U$$4156/B1 U$$4182/B2 VGND VGND VPWR VPWR U$$4157/A sky130_fd_sc_hd__a22o_1
XFILLER_24_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3411 U$$3411/A U$$3423/B VGND VGND VPWR VPWR U$$3411/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_113_1 input144/X dadda_fa_4_113_1/B dadda_fa_4_113_1/CIN VGND VGND VPWR
+ VPWR dadda_fa_5_114_0/B dadda_fa_5_113_1/B sky130_fd_sc_hd__fa_1
XU$$3422 U$$4516/B1 U$$3292/X U$$3422/B1 U$$3293/X VGND VGND VPWR VPWR U$$3423/A sky130_fd_sc_hd__a22o_1
XFILLER_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4167 U$$4167/A U$$4215/B VGND VGND VPWR VPWR U$$4167/X sky130_fd_sc_hd__xor2_1
XU$$3433 U$$3844/A1 U$$3479/A2 U$$3709/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3434/A
+ sky130_fd_sc_hd__a22o_1
XU$$4178 _582_/Q U$$4202/A2 U$$4180/A1 U$$4202/B2 VGND VGND VPWR VPWR U$$4179/A sky130_fd_sc_hd__a22o_1
XU$$4189 U$$4189/A U$$4197/B VGND VGND VPWR VPWR U$$4189/X sky130_fd_sc_hd__xor2_1
XU$$3444 U$$3444/A U$$3478/B VGND VGND VPWR VPWR U$$3444/X sky130_fd_sc_hd__xor2_1
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3455 U$$4003/A1 U$$3559/A2 U$$4140/B1 U$$3559/B2 VGND VGND VPWR VPWR U$$3456/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2710 U$$2710/A U$$2739/A VGND VGND VPWR VPWR U$$2710/X sky130_fd_sc_hd__xor2_1
XU$$2721 U$$2858/A1 U$$2729/A2 U$$2721/B1 U$$2729/B2 VGND VGND VPWR VPWR U$$2722/A
+ sky130_fd_sc_hd__a22o_1
XU$$3466 U$$3466/A U$$3561/A VGND VGND VPWR VPWR U$$3466/X sky130_fd_sc_hd__xor2_1
XFILLER_80_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_106_0 dadda_fa_4_106_0/A dadda_fa_4_106_0/B dadda_fa_4_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/A dadda_fa_5_106_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_39_5 dadda_fa_2_39_5/A dadda_fa_2_39_5/B dadda_fa_2_39_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_40_2/A dadda_fa_4_39_0/A sky130_fd_sc_hd__fa_2
XU$$2732 U$$2732/A U$$2734/B VGND VGND VPWR VPWR U$$2732/X sky130_fd_sc_hd__xor2_1
XFILLER_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3477 U$$4160/B1 U$$3479/A2 U$$4027/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3478/A
+ sky130_fd_sc_hd__a22o_1
XU$$3488 U$$3488/A U$$3520/B VGND VGND VPWR VPWR U$$3488/X sky130_fd_sc_hd__xor2_1
XFILLER_18_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2743 U$$2877/A U$$2743/B VGND VGND VPWR VPWR U$$2743/X sky130_fd_sc_hd__and2_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2754 U$$2754/A1 U$$2788/A2 U$$2756/A1 U$$2788/B2 VGND VGND VPWR VPWR U$$2755/A
+ sky130_fd_sc_hd__a22o_1
XU$$3499 U$$3771/B1 U$$3545/A2 U$$3638/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3500/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2765 U$$2765/A U$$2813/B VGND VGND VPWR VPWR U$$2765/X sky130_fd_sc_hd__xor2_1
XFILLER_61_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2776 U$$4418/B1 U$$2814/A2 U$$4285/A1 U$$2814/B2 VGND VGND VPWR VPWR U$$2777/A
+ sky130_fd_sc_hd__a22o_1
XU$$2787 U$$2787/A U$$2787/B VGND VGND VPWR VPWR U$$2787/X sky130_fd_sc_hd__xor2_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2798 U$$4305/A1 U$$2798/A2 U$$4168/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2799/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_99_1 dadda_fa_5_99_1/A dadda_fa_5_99_1/B dadda_fa_5_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_100_0/B dadda_fa_7_99_0/A sky130_fd_sc_hd__fa_1
XFILLER_190_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_894 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4451_1804 VGND VGND VPWR VPWR U$$4451_1804/HI U$$4451/B sky130_fd_sc_hd__conb_1
XFILLER_142_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$705 final_adder.U$$705/A final_adder.U$$705/B VGND VGND VPWR VPWR
+ _251_/D sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$716 final_adder.U$$716/A final_adder.U$$716/B VGND VGND VPWR VPWR
+ _262_/D sky130_fd_sc_hd__xor2_1
XFILLER_84_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater920 _677_/Q VGND VGND VPWR VPWR U$$4203/B sky130_fd_sc_hd__buf_4
XFILLER_112_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$727 final_adder.U$$727/A final_adder.U$$727/B VGND VGND VPWR VPWR
+ _273_/D sky130_fd_sc_hd__xor2_4
Xrepeater931 U$$3895/B VGND VGND VPWR VPWR U$$3873/B sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$738 final_adder.U$$738/A final_adder.U$$738/B VGND VGND VPWR VPWR
+ _284_/D sky130_fd_sc_hd__xor2_4
XFILLER_111_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater942 U$$3804/B VGND VGND VPWR VPWR U$$3800/B sky130_fd_sc_hd__buf_8
XFILLER_56_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$749 final_adder.U$$749/A final_adder.U$$749/B VGND VGND VPWR VPWR
+ _295_/D sky130_fd_sc_hd__xor2_4
XFILLER_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater953 _669_/Q VGND VGND VPWR VPWR U$$3699/A sky130_fd_sc_hd__buf_6
XFILLER_99_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater964 U$$3562/A VGND VGND VPWR VPWR U$$3538/B sky130_fd_sc_hd__buf_6
XFILLER_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater975 U$$3276/B VGND VGND VPWR VPWR U$$3232/B sky130_fd_sc_hd__buf_8
Xrepeater986 U$$3077/B VGND VGND VPWR VPWR U$$3083/B sky130_fd_sc_hd__buf_6
XFILLER_204_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater997 U$$3008/B VGND VGND VPWR VPWR U$$3000/B sky130_fd_sc_hd__buf_8
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_583 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_439 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_94_0 dadda_fa_4_94_0/A dadda_fa_4_94_0/B dadda_fa_4_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/A dadda_fa_5_94_1/A sky130_fd_sc_hd__fa_1
XFILLER_119_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_108_2 U$$4080/X U$$4213/X U$$4346/X VGND VGND VPWR VPWR dadda_fa_4_109_1/A
+ dadda_fa_4_108_2/B sky130_fd_sc_hd__fa_1
XFILLER_106_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput280 _288_/Q VGND VGND VPWR VPWR o[120] sky130_fd_sc_hd__buf_2
XFILLER_0_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput291 _183_/Q VGND VGND VPWR VPWR o[15] sky130_fd_sc_hd__buf_2
XFILLER_43_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2006 U$$2963/B1 U$$2040/A2 U$$4474/A1 U$$2040/B2 VGND VGND VPWR VPWR U$$2007/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2017 U$$2017/A U$$2029/B VGND VGND VPWR VPWR U$$2017/X sky130_fd_sc_hd__xor2_1
XU$$2028 U$$382/B1 U$$2028/A2 U$$384/B1 U$$2028/B2 VGND VGND VPWR VPWR U$$2029/A sky130_fd_sc_hd__a22o_1
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2039 U$$2039/A U$$2039/B VGND VGND VPWR VPWR U$$2039/X sky130_fd_sc_hd__xor2_1
XFILLER_204_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1305 U$$3221/B1 U$$1309/A2 U$$3088/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1306/A
+ sky130_fd_sc_hd__a22o_1
XU$$1316 U$$1316/A U$$1356/B VGND VGND VPWR VPWR U$$1316/X sky130_fd_sc_hd__xor2_1
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1327 U$$94/A1 U$$1237/X U$$2971/B1 U$$1238/X VGND VGND VPWR VPWR U$$1328/A sky130_fd_sc_hd__a22o_1
XFILLER_167_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1338 U$$1338/A U$$1370/A VGND VGND VPWR VPWR U$$1338/X sky130_fd_sc_hd__xor2_1
XU$$1349 U$$527/A1 U$$1367/A2 U$$253/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1350/A sky130_fd_sc_hd__a22o_1
XFILLER_128_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_731 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_206_ _213_/CLK _206_/D VGND VGND VPWR VPWR _206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_51_4 dadda_fa_2_51_4/A dadda_fa_2_51_4/B dadda_fa_2_51_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/CIN dadda_fa_3_51_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_44_3 dadda_fa_2_44_3/A dadda_fa_2_44_3/B dadda_fa_2_44_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_1/B dadda_fa_3_44_3/B sky130_fd_sc_hd__fa_1
XFILLER_65_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3230 U$$3230/A U$$3232/B VGND VGND VPWR VPWR U$$3230/X sky130_fd_sc_hd__xor2_1
XFILLER_19_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$12 _436_/Q _308_/Q VGND VGND VPWR VPWR final_adder.U$$507/B1 final_adder.U$$634/A
+ sky130_fd_sc_hd__ha_2
XU$$3241 U$$4474/A1 U$$3283/A2 U$$4476/A1 U$$3283/B2 VGND VGND VPWR VPWR U$$3242/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_640 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$23 _447_/Q _319_/Q VGND VGND VPWR VPWR final_adder.U$$151/B1 final_adder.U$$645/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$34 _458_/Q _330_/Q VGND VGND VPWR VPWR final_adder.U$$529/B1 final_adder.U$$656/A
+ sky130_fd_sc_hd__ha_1
XU$$3252 U$$3252/A U$$3256/B VGND VGND VPWR VPWR U$$3252/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_37_2 U$$1544/X U$$1677/X U$$1810/X VGND VGND VPWR VPWR dadda_fa_3_38_1/A
+ dadda_fa_3_37_3/A sky130_fd_sc_hd__fa_1
XU$$4481_1819 VGND VGND VPWR VPWR U$$4481_1819/HI U$$4481/B sky130_fd_sc_hd__conb_1
XFILLER_65_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3263 _604_/Q U$$3263/A2 U$$3539/A1 U$$3263/B2 VGND VGND VPWR VPWR U$$3264/A sky130_fd_sc_hd__a22o_1
XFILLER_81_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$45 _469_/Q _341_/Q VGND VGND VPWR VPWR final_adder.U$$173/B1 final_adder.U$$667/A
+ sky130_fd_sc_hd__ha_2
XU$$3274 U$$3274/A U$$3276/B VGND VGND VPWR VPWR U$$3274/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$56 _480_/Q _352_/Q VGND VGND VPWR VPWR final_adder.U$$551/B1 final_adder.U$$678/A
+ sky130_fd_sc_hd__ha_1
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3285 U$$3285/A1 U$$3285/A2 U$$3285/B1 U$$3285/B2 VGND VGND VPWR VPWR U$$3286/A
+ sky130_fd_sc_hd__a22o_1
XU$$2540 U$$3362/A1 U$$2566/A2 U$$3362/B1 U$$2566/B2 VGND VGND VPWR VPWR U$$2541/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2551 U$$2551/A U$$2551/B VGND VGND VPWR VPWR U$$2551/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_14_1 dadda_fa_5_14_1/A dadda_fa_5_14_1/B dadda_fa_5_14_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_15_0/B dadda_fa_7_14_0/A sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$67 _491_/Q _363_/Q VGND VGND VPWR VPWR final_adder.U$$195/B1 final_adder.U$$689/A
+ sky130_fd_sc_hd__ha_2
XFILLER_94_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$78 _502_/Q _374_/Q VGND VGND VPWR VPWR final_adder.U$$573/B1 final_adder.U$$700/A
+ sky130_fd_sc_hd__ha_1
XFILLER_146_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3296 _552_/Q U$$3320/A2 U$$3709/A1 U$$3320/B2 VGND VGND VPWR VPWR U$$3297/A sky130_fd_sc_hd__a22o_1
XFILLER_185_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2562 U$$3932/A1 U$$2588/A2 U$$918/B1 U$$2588/B2 VGND VGND VPWR VPWR U$$2563/A
+ sky130_fd_sc_hd__a22o_1
XU$$2573 U$$2573/A U$$2583/B VGND VGND VPWR VPWR U$$2573/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$89 _513_/Q _385_/Q VGND VGND VPWR VPWR final_adder.U$$217/B1 final_adder.U$$711/A
+ sky130_fd_sc_hd__ha_2
XU$$2584 U$$3132/A1 U$$2588/A2 U$$3132/B1 U$$2588/B2 VGND VGND VPWR VPWR U$$2585/A
+ sky130_fd_sc_hd__a22o_1
XU$$4409_1783 VGND VGND VPWR VPWR U$$4409_1783/HI U$$4409/B sky130_fd_sc_hd__conb_1
XU$$2595 U$$2595/A U$$2597/B VGND VGND VPWR VPWR U$$2595/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1850 U$$1850/A U$$1852/B VGND VGND VPWR VPWR U$$1850/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1861 U$$491/A1 U$$1785/X U$$493/A1 U$$1786/X VGND VGND VPWR VPWR U$$1862/A sky130_fd_sc_hd__a22o_1
XFILLER_179_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1872 U$$1872/A U$$1918/A VGND VGND VPWR VPWR U$$1872/X sky130_fd_sc_hd__xor2_1
XFILLER_107_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1883 U$$3388/B1 U$$1915/A2 U$$3253/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1884/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1894 U$$1894/A U$$1917/A VGND VGND VPWR VPWR U$$1894/X sky130_fd_sc_hd__xor2_1
XFILLER_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_945 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1110 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$513 final_adder.U$$640/A final_adder.U$$640/B final_adder.U$$513/B1
+ VGND VGND VPWR VPWR final_adder.U$$641/B sky130_fd_sc_hd__a21o_1
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$535 final_adder.U$$662/A final_adder.U$$662/B final_adder.U$$535/B1
+ VGND VGND VPWR VPWR final_adder.U$$663/B sky130_fd_sc_hd__a21o_1
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater750 U$$3066/B2 VGND VGND VPWR VPWR U$$3054/B2 sky130_fd_sc_hd__buf_4
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$557 final_adder.U$$684/A final_adder.U$$684/B final_adder.U$$557/B1
+ VGND VGND VPWR VPWR final_adder.U$$685/B sky130_fd_sc_hd__a21o_1
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater761 U$$2981/B2 VGND VGND VPWR VPWR U$$2943/B2 sky130_fd_sc_hd__buf_6
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$407 U$$407/A _621_/Q VGND VGND VPWR VPWR U$$407/X sky130_fd_sc_hd__xor2_1
Xrepeater772 U$$392/B2 VGND VGND VPWR VPWR U$$384/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$579 final_adder.U$$706/A final_adder.U$$706/B final_adder.U$$579/B1
+ VGND VGND VPWR VPWR final_adder.U$$707/B sky130_fd_sc_hd__a21o_1
XU$$418 U$$418/A U$$452/B VGND VGND VPWR VPWR U$$418/X sky130_fd_sc_hd__xor2_1
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater783 U$$2707/B2 VGND VGND VPWR VPWR U$$2697/B2 sky130_fd_sc_hd__buf_6
Xrepeater794 U$$2530/B2 VGND VGND VPWR VPWR U$$2524/B2 sky130_fd_sc_hd__buf_4
XU$$429 U$$429/A1 U$$457/A2 U$$429/B1 U$$457/B2 VGND VGND VPWR VPWR U$$430/A sky130_fd_sc_hd__a22o_1
XFILLER_204_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1307 U$$3255/B1 VGND VGND VPWR VPWR U$$791/A1 sky130_fd_sc_hd__buf_6
XFILLER_197_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_113_0 U$$3424/Y U$$3558/X U$$3691/X VGND VGND VPWR VPWR dadda_fa_4_114_1/CIN
+ dadda_fa_4_113_2/B sky130_fd_sc_hd__fa_1
XFILLER_181_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1318 U$$4214/A1 VGND VGND VPWR VPWR U$$926/A1 sky130_fd_sc_hd__buf_6
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1329 U$$4075/A1 VGND VGND VPWR VPWR U$$4486/A1 sky130_fd_sc_hd__buf_6
XFILLER_69_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_61_3 dadda_fa_3_61_3/A dadda_fa_3_61_3/B dadda_fa_3_61_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_1/B dadda_fa_4_61_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_94_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_54_2 dadda_fa_3_54_2/A dadda_fa_3_54_2/B dadda_fa_3_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_1/A dadda_fa_4_54_2/B sky130_fd_sc_hd__fa_1
XFILLER_134_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_47_1 dadda_fa_3_47_1/A dadda_fa_3_47_1/B dadda_fa_3_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_0/CIN dadda_fa_4_47_2/A sky130_fd_sc_hd__fa_1
XFILLER_75_475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_24_0 dadda_fa_6_24_0/A dadda_fa_6_24_0/B dadda_fa_6_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_25_0/B dadda_fa_7_24_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_870 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$930 U$$930/A1 U$$826/X U$$932/A1 U$$827/X VGND VGND VPWR VPWR U$$931/A sky130_fd_sc_hd__a22o_1
XU$$941 U$$941/A U$$951/B VGND VGND VPWR VPWR U$$941/X sky130_fd_sc_hd__xor2_1
XFILLER_211_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$952 U$$952/A1 U$$956/A2 U$$954/A1 U$$956/B2 VGND VGND VPWR VPWR U$$953/A sky130_fd_sc_hd__a22o_1
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$963 U$$961/Y _630_/Q _629_/Q U$$962/X U$$959/Y VGND VGND VPWR VPWR U$$963/X sky130_fd_sc_hd__a32o_4
XU$$1102 U$$1102/A1 U$$1194/A2 U$$967/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1103/A
+ sky130_fd_sc_hd__a22o_1
XU$$1113 U$$1113/A U$$1147/B VGND VGND VPWR VPWR U$$1113/X sky130_fd_sc_hd__xor2_1
XU$$974 U$$974/A U$$994/B VGND VGND VPWR VPWR U$$974/X sky130_fd_sc_hd__xor2_1
XU$$1124 U$$302/A1 U$$1150/A2 U$$989/A1 U$$1150/B2 VGND VGND VPWR VPWR U$$1125/A sky130_fd_sc_hd__a22o_1
XFILLER_16_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$985 U$$985/A1 U$$997/A2 U$$987/A1 U$$997/B2 VGND VGND VPWR VPWR U$$986/A sky130_fd_sc_hd__a22o_1
XU$$1135 U$$1135/A U$$1147/B VGND VGND VPWR VPWR U$$1135/X sky130_fd_sc_hd__xor2_1
XU$$996 U$$996/A U$$996/B VGND VGND VPWR VPWR U$$996/X sky130_fd_sc_hd__xor2_1
XFILLER_44_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1006 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1146 U$$48/B1 U$$1146/A2 U$$874/A1 U$$1146/B2 VGND VGND VPWR VPWR U$$1147/A sky130_fd_sc_hd__a22o_1
XFILLER_44_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1157 U$$1157/A U$$1191/B VGND VGND VPWR VPWR U$$1157/X sky130_fd_sc_hd__xor2_1
XU$$1168 U$$72/A1 U$$1176/A2 U$$74/A1 U$$1176/B2 VGND VGND VPWR VPWR U$$1169/A sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_112_2 U$$4088/X U$$4221/X VGND VGND VPWR VPWR dadda_fa_4_113_2/A dadda_ha_3_112_2/SUM
+ sky130_fd_sc_hd__ha_1
XU$$1179 U$$1179/A U$$1225/B VGND VGND VPWR VPWR U$$1179/X sky130_fd_sc_hd__xor2_1
XFILLER_176_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_580 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_639 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_99_4 U$$4062/X U$$4195/X U$$4328/X VGND VGND VPWR VPWR dadda_fa_3_100_2/B
+ dadda_fa_4_99_0/A sky130_fd_sc_hd__fa_1
XFILLER_160_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4439_1798 VGND VGND VPWR VPWR U$$4439_1798/HI U$$4439/B sky130_fd_sc_hd__conb_1
XFILLER_171_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_42_0 U$$1953/X U$$2086/X U$$2219/X VGND VGND VPWR VPWR dadda_fa_3_43_0/B
+ dadda_fa_3_42_2/B sky130_fd_sc_hd__fa_1
XFILLER_54_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3060 U$$4430/A1 U$$3066/A2 U$$4432/A1 U$$3066/B2 VGND VGND VPWR VPWR U$$3061/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3071 U$$3071/A U$$3107/B VGND VGND VPWR VPWR U$$3071/X sky130_fd_sc_hd__xor2_1
XU$$3082 U$$3354/B1 U$$3082/A2 U$$3221/A1 U$$3082/B2 VGND VGND VPWR VPWR U$$3083/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3093 U$$3093/A U$$3121/B VGND VGND VPWR VPWR U$$3093/X sky130_fd_sc_hd__xor2_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2370 U$$2370/A U$$2418/B VGND VGND VPWR VPWR U$$2370/X sky130_fd_sc_hd__xor2_1
XFILLER_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_5__f_clk clkbuf_2_2_0_clk/X VGND VGND VPWR VPWR _628_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2381 U$$3475/B1 U$$2387/A2 U$$3342/A1 U$$2387/B2 VGND VGND VPWR VPWR U$$2382/A
+ sky130_fd_sc_hd__a22o_1
XU$$2392 U$$2392/A U$$2400/B VGND VGND VPWR VPWR U$$2392/X sky130_fd_sc_hd__xor2_1
XFILLER_210_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1680 U$$310/A1 U$$1740/A2 U$$584/B1 U$$1740/B2 VGND VGND VPWR VPWR U$$1681/A sky130_fd_sc_hd__a22o_1
XFILLER_14_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1691 U$$1691/A U$$1723/B VGND VGND VPWR VPWR U$$1691/X sky130_fd_sc_hd__xor2_1
XFILLER_194_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_88_4 U$$3242/X U$$3375/X VGND VGND VPWR VPWR dadda_fa_2_89_4/CIN dadda_fa_3_88_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_148_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_71_2 dadda_fa_4_71_2/A dadda_fa_4_71_2/B dadda_fa_4_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/CIN dadda_fa_5_71_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_87_2 U$$2442/X U$$2575/X U$$2708/X VGND VGND VPWR VPWR dadda_fa_2_88_3/CIN
+ dadda_fa_2_87_5/B sky130_fd_sc_hd__fa_1
XFILLER_39_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_64_1 dadda_fa_4_64_1/A dadda_fa_4_64_1/B dadda_fa_4_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/B dadda_fa_5_64_1/B sky130_fd_sc_hd__fa_1
XFILLER_89_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_41_0 dadda_fa_7_41_0/A dadda_fa_7_41_0/B dadda_fa_7_41_0/CIN VGND VGND
+ VPWR VPWR _466_/D _337_/D sky130_fd_sc_hd__fa_1
XFILLER_77_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_57_0 dadda_fa_4_57_0/A dadda_fa_4_57_0/B dadda_fa_4_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/A dadda_fa_5_57_1/A sky130_fd_sc_hd__fa_1
XFILLER_44_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_420 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$310 final_adder.U$$310/A final_adder.U$$310/B VGND VGND VPWR VPWR
+ final_adder.U$$346/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$321 final_adder.U$$258/X final_adder.U$$626/B final_adder.U$$259/X
+ VGND VGND VPWR VPWR final_adder.U$$630/B sky130_fd_sc_hd__a21o_4
XFILLER_131_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$332 final_adder.U$$332/A final_adder.U$$332/B VGND VGND VPWR VPWR
+ final_adder.U$$358/B sky130_fd_sc_hd__and2_1
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$343 final_adder.U$$342/A final_adder.U$$301/X final_adder.U$$303/X
+ VGND VGND VPWR VPWR final_adder.U$$343/X sky130_fd_sc_hd__a21o_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$354 final_adder.U$$354/A final_adder.U$$354/B VGND VGND VPWR VPWR
+ final_adder.U$$354/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$365 final_adder.U$$364/A final_adder.U$$345/X ANTENNA_10/DIODE VGND
+ VGND VPWR VPWR final_adder.U$$365/X sky130_fd_sc_hd__a21o_1
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$204 U$$204/A U$$216/B VGND VGND VPWR VPWR U$$204/X sky130_fd_sc_hd__xor2_1
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater580 U$$2040/A2 VGND VGND VPWR VPWR U$$2038/A2 sky130_fd_sc_hd__buf_6
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$215 U$$900/A1 U$$217/A2 U$$80/A1 U$$217/B2 VGND VGND VPWR VPWR U$$216/A sky130_fd_sc_hd__a22o_1
X_540_ _541_/CLK _540_/D VGND VGND VPWR VPWR _540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$387 final_adder.U$$372/B final_adder.U$$686/B final_adder.U$$361/X
+ VGND VGND VPWR VPWR final_adder.U$$702/B sky130_fd_sc_hd__a21o_1
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater591 U$$1736/A2 VGND VGND VPWR VPWR U$$1684/A2 sky130_fd_sc_hd__buf_4
XU$$226 U$$226/A U$$226/B VGND VGND VPWR VPWR U$$226/X sky130_fd_sc_hd__xor2_1
XFILLER_45_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$237 U$$648/A1 U$$249/A2 U$$648/B1 U$$249/B2 VGND VGND VPWR VPWR U$$238/A sky130_fd_sc_hd__a22o_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$248 U$$248/A U$$250/B VGND VGND VPWR VPWR U$$248/X sky130_fd_sc_hd__xor2_1
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$259 U$$942/B1 U$$259/A2 U$$946/A1 U$$259/B2 VGND VGND VPWR VPWR U$$260/A sky130_fd_sc_hd__a22o_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_471_ _471_/CLK _471_/D VGND VGND VPWR VPWR _471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1083 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_303 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$9 U$$9/A U$$9/B VGND VGND VPWR VPWR U$$9/X sky130_fd_sc_hd__xor2_1
XFILLER_138_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1104 U$$1296/B VGND VGND VPWR VPWR U$$1310/B sky130_fd_sc_hd__buf_6
XFILLER_126_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1115 U$$1203/B VGND VGND VPWR VPWR U$$1195/B sky130_fd_sc_hd__buf_6
Xrepeater1126 U$$1095/A VGND VGND VPWR VPWR U$$1090/B sky130_fd_sc_hd__buf_6
Xrepeater1137 _629_/Q VGND VGND VPWR VPWR U$$935/B sky130_fd_sc_hd__buf_8
Xrepeater1148 U$$684/A VGND VGND VPWR VPWR U$$651/B sky130_fd_sc_hd__buf_6
Xrepeater1159 U$$536/B VGND VGND VPWR VPWR U$$500/B sky130_fd_sc_hd__buf_6
XFILLER_101_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_102_0_1863 VGND VGND VPWR VPWR dadda_fa_2_102_0/A dadda_fa_2_102_0_1863/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_106_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_75_0 U$$821/Y U$$955/X U$$1088/X VGND VGND VPWR VPWR dadda_fa_1_76_8/A
+ dadda_fa_1_75_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$760 U$$760/A U$$760/B VGND VGND VPWR VPWR U$$760/X sky130_fd_sc_hd__xor2_1
XFILLER_90_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_669_ _674_/CLK _669_/D VGND VGND VPWR VPWR _669_/Q sky130_fd_sc_hd__dfxtp_4
XU$$771 U$$84/B1 U$$783/A2 U$$910/A1 U$$783/B2 VGND VGND VPWR VPWR U$$772/A sky130_fd_sc_hd__a22o_1
XFILLER_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$782 U$$782/A U$$821/A VGND VGND VPWR VPWR U$$782/X sky130_fd_sc_hd__xor2_1
XU$$793 U$$930/A1 U$$795/A2 U$$932/A1 U$$795/B2 VGND VGND VPWR VPWR U$$794/A sky130_fd_sc_hd__a22o_1
XFILLER_50_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_81_1 dadda_fa_5_81_1/A dadda_fa_5_81_1/B dadda_fa_5_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_82_0/B dadda_fa_7_81_0/A sky130_fd_sc_hd__fa_2
XFILLER_117_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_97_1 U$$2728/X U$$2861/X U$$2994/X VGND VGND VPWR VPWR dadda_fa_3_98_0/CIN
+ dadda_fa_3_97_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_74_0 dadda_fa_5_74_0/A dadda_fa_5_74_0/B dadda_fa_5_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_75_0/A dadda_fa_6_74_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1660 U$$4404/A1 VGND VGND VPWR VPWR U$$3445/A1 sky130_fd_sc_hd__buf_6
XFILLER_104_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1671 U$$2345/A1 VGND VGND VPWR VPWR U$$16/A1 sky130_fd_sc_hd__buf_6
Xrepeater1682 U$$3163/B1 VGND VGND VPWR VPWR U$$2754/A1 sky130_fd_sc_hd__buf_4
XFILLER_116_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1693 U$$3437/A1 VGND VGND VPWR VPWR U$$3024/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_73_8 dadda_fa_1_73_8/A dadda_fa_1_73_8/B dadda_fa_1_73_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_74_3/A dadda_fa_3_73_0/A sky130_fd_sc_hd__fa_2
XFILLER_59_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_494 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_66_7 dadda_fa_1_66_7/A dadda_fa_1_66_7/B dadda_fa_1_66_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_2/CIN dadda_fa_2_66_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_59_6 U$$3982/X input211/X dadda_fa_1_59_6/CIN VGND VGND VPWR VPWR dadda_fa_2_60_2/B
+ dadda_fa_2_59_5/B sky130_fd_sc_hd__fa_1
XFILLER_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_89_0 dadda_fa_7_89_0/A dadda_fa_7_89_0/B dadda_fa_7_89_0/CIN VGND VGND
+ VPWR VPWR _514_/D _385_/D sky130_fd_sc_hd__fa_1
XFILLER_175_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_92_0 dadda_fa_1_92_0/A U$$2053/X U$$2186/X VGND VGND VPWR VPWR dadda_fa_2_93_4/CIN
+ dadda_fa_2_92_5/B sky130_fd_sc_hd__fa_1
XFILLER_11_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4508 U$$4508/A1 U$$4388/X U$$4510/A1 U$$4516/B2 VGND VGND VPWR VPWR U$$4509/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$140 final_adder.U$$635/A final_adder.U$$634/A VGND VGND VPWR VPWR
+ final_adder.U$$262/B sky130_fd_sc_hd__and2_1
XU$$3807 U$$4218/A1 U$$3823/A2 U$$3807/B1 U$$3823/B2 VGND VGND VPWR VPWR U$$3808/A
+ sky130_fd_sc_hd__a22o_1
XU$$3818 U$$3818/A U$$3835/A VGND VGND VPWR VPWR U$$3818/X sky130_fd_sc_hd__xor2_1
XFILLER_57_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3829 U$$4238/B1 U$$3833/A2 U$$406/A1 U$$3833/B2 VGND VGND VPWR VPWR U$$3830/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$151 final_adder.U$$645/A final_adder.U$$517/B1 final_adder.U$$151/B1
+ VGND VGND VPWR VPWR final_adder.U$$151/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$162 final_adder.U$$657/A final_adder.U$$656/A VGND VGND VPWR VPWR
+ final_adder.U$$272/A sky130_fd_sc_hd__and2_1
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_104_0 dadda_fa_6_104_0/A dadda_fa_6_104_0/B dadda_fa_6_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_105_0/B dadda_fa_7_104_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$173 final_adder.U$$667/A final_adder.U$$539/B1 final_adder.U$$173/B1
+ VGND VGND VPWR VPWR final_adder.U$$173/X sky130_fd_sc_hd__a21o_1
XFILLER_85_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$184 final_adder.U$$679/A final_adder.U$$678/A VGND VGND VPWR VPWR
+ final_adder.U$$284/B sky130_fd_sc_hd__and2_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$195 final_adder.U$$689/A final_adder.U$$561/B1 final_adder.U$$195/B1
+ VGND VGND VPWR VPWR final_adder.U$$195/X sky130_fd_sc_hd__a21o_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_523_ _523_/CLK _523_/D VGND VGND VPWR VPWR _523_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_24_3 input173/X dadda_fa_3_24_3/B dadda_fa_3_24_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_25_1/B dadda_fa_4_24_2/CIN sky130_fd_sc_hd__fa_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_454_ _454_/CLK _454_/D VGND VGND VPWR VPWR _454_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_385_ _515_/CLK _385_/D VGND VGND VPWR VPWR _385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_91_0 dadda_fa_6_91_0/A dadda_fa_6_91_0/B dadda_fa_6_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_92_0/B dadda_fa_7_91_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_103_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_835 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_69_5 dadda_fa_2_69_5/A dadda_fa_2_69_5/B dadda_fa_2_69_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_2/A dadda_fa_4_69_0/A sky130_fd_sc_hd__fa_1
XFILLER_114_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput180 c[30] VGND VGND VPWR VPWR input180/X sky130_fd_sc_hd__clkbuf_1
Xinput191 c[40] VGND VGND VPWR VPWR input191/X sky130_fd_sc_hd__buf_2
XFILLER_48_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$590 U$$42/A1 U$$622/A2 U$$42/B1 U$$622/B2 VGND VGND VPWR VPWR U$$591/A sky130_fd_sc_hd__a22o_1
XFILLER_211_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_194 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_390 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1490 U$$3624/A1 VGND VGND VPWR VPWR U$$4444/B1 sky130_fd_sc_hd__buf_8
XFILLER_28_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_71_5 U$$4139/X U$$4272/X U$$4405/X VGND VGND VPWR VPWR dadda_fa_2_72_2/A
+ dadda_fa_2_71_5/A sky130_fd_sc_hd__fa_1
XFILLER_101_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_64_4 U$$4125/X U$$4258/X U$$4391/X VGND VGND VPWR VPWR dadda_fa_2_65_1/CIN
+ dadda_fa_2_64_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_57_3 U$$2382/X U$$2515/X U$$2648/X VGND VGND VPWR VPWR dadda_fa_2_58_1/B
+ dadda_fa_2_57_4/B sky130_fd_sc_hd__fa_1
XFILLER_27_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_34_2 dadda_fa_4_34_2/A dadda_fa_4_34_2/B dadda_fa_4_34_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/CIN dadda_fa_5_34_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_27_1 dadda_fa_4_27_1/A dadda_fa_4_27_1/B dadda_fa_4_27_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/B dadda_fa_5_27_1/B sky130_fd_sc_hd__fa_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ _179_/CLK _170_/D VGND VGND VPWR VPWR _170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4305 U$$4305/A1 U$$4347/A2 U$$4444/A1 U$$4347/B2 VGND VGND VPWR VPWR U$$4306/A
+ sky130_fd_sc_hd__a22o_1
XU$$4316 U$$4316/A U$$4322/B VGND VGND VPWR VPWR U$$4316/X sky130_fd_sc_hd__xor2_1
XFILLER_120_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4327 U$$4464/A1 U$$4327/A2 U$$4466/A1 U$$4333/B2 VGND VGND VPWR VPWR U$$4328/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4338 U$$4338/A U$$4350/B VGND VGND VPWR VPWR U$$4338/X sky130_fd_sc_hd__xor2_1
XFILLER_93_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4349 U$$4486/A1 U$$4381/A2 U$$4351/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4350/A
+ sky130_fd_sc_hd__a22o_1
XU$$3604 U$$3876/B1 U$$3628/A2 U$$4291/A1 U$$3628/B2 VGND VGND VPWR VPWR U$$3605/A
+ sky130_fd_sc_hd__a22o_1
XU$$3615 U$$3615/A U$$3627/B VGND VGND VPWR VPWR U$$3615/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_16_1 U$$438/X U$$571/X VGND VGND VPWR VPWR dadda_fa_4_17_2/A dadda_ha_3_16_1/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3626 U$$4448/A1 U$$3662/A2 U$$3626/B1 U$$3662/B2 VGND VGND VPWR VPWR U$$3627/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3637 U$$3637/A U$$3637/B VGND VGND VPWR VPWR U$$3637/X sky130_fd_sc_hd__xor2_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2903 U$$4410/A1 U$$2959/A2 U$$3042/A1 U$$2959/B2 VGND VGND VPWR VPWR U$$2904/A
+ sky130_fd_sc_hd__a22o_1
XU$$3648 U$$4194/B1 U$$3662/A2 U$$4061/A1 U$$3662/B2 VGND VGND VPWR VPWR U$$3649/A
+ sky130_fd_sc_hd__a22o_1
XU$$3659 U$$3659/A U$$3671/B VGND VGND VPWR VPWR U$$3659/X sky130_fd_sc_hd__xor2_1
XU$$2914 U$$2914/A U$$2916/B VGND VGND VPWR VPWR U$$2914/X sky130_fd_sc_hd__xor2_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2925 U$$596/A1 U$$2929/A2 U$$596/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2926/A sky130_fd_sc_hd__a22o_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2936 U$$2936/A U$$2972/B VGND VGND VPWR VPWR U$$2936/X sky130_fd_sc_hd__xor2_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2947 U$$3358/A1 U$$2981/A2 U$$2947/B1 U$$2981/B2 VGND VGND VPWR VPWR U$$2948/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_230 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_22_0 U$$317/X U$$450/X U$$583/X VGND VGND VPWR VPWR dadda_fa_4_23_0/B
+ dadda_fa_4_22_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_209_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2958 U$$2958/A U$$2982/B VGND VGND VPWR VPWR U$$2958/X sky130_fd_sc_hd__xor2_1
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_241 _192_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_506_ _507_/CLK _506_/D VGND VGND VPWR VPWR _506_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2969 U$$4476/A1 U$$2973/A2 U$$4478/A1 U$$2973/B2 VGND VGND VPWR VPWR U$$2970/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_252 _195_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_263 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 _212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 _214_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_296 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_437_ _444_/CLK _437_/D VGND VGND VPWR VPWR _437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_368_ _634_/CLK _368_/D VGND VGND VPWR VPWR _368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_299_ _428_/CLK _299_/D VGND VGND VPWR VPWR _299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_832 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_81_4 dadda_fa_2_81_4/A dadda_fa_2_81_4/B dadda_fa_2_81_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/CIN dadda_fa_3_81_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_74_3 dadda_fa_2_74_3/A dadda_fa_2_74_3/B dadda_fa_2_74_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/B dadda_fa_3_74_3/B sky130_fd_sc_hd__fa_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_67_2 dadda_fa_2_67_2/A dadda_fa_2_67_2/B dadda_fa_2_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/A dadda_fa_3_67_3/A sky130_fd_sc_hd__fa_1
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_44_1 dadda_fa_5_44_1/A dadda_fa_5_44_1/B dadda_fa_5_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_45_0/B dadda_fa_7_44_0/A sky130_fd_sc_hd__fa_1
XFILLER_28_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_37_0 dadda_fa_5_37_0/A dadda_fa_5_37_0/B dadda_fa_5_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_38_0/A dadda_fa_6_37_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_111_0 dadda_fa_5_111_0/A dadda_fa_5_111_0/B dadda_fa_5_111_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_112_0/A dadda_fa_6_111_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_1 U$$2791/X U$$2924/X U$$3057/X VGND VGND VPWR VPWR dadda_fa_2_63_0/CIN
+ dadda_fa_2_62_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_41_1030 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_55_0 U$$782/X U$$915/X U$$1048/X VGND VGND VPWR VPWR dadda_fa_2_56_0/B
+ dadda_fa_2_55_3/B sky130_fd_sc_hd__fa_1
XFILLER_86_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1509 U$$1642/B VGND VGND VPWR VPWR U$$1509/Y sky130_fd_sc_hd__inv_1
XFILLER_203_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_222_ _225_/CLK _222_/D VGND VGND VPWR VPWR _222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_91_3 dadda_fa_3_91_3/A dadda_fa_3_91_3/B dadda_fa_3_91_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_1/B dadda_fa_4_91_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_183_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_84_2 dadda_fa_3_84_2/A dadda_fa_3_84_2/B dadda_fa_3_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_1/A dadda_fa_4_84_2/B sky130_fd_sc_hd__fa_1
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_77_1 dadda_fa_3_77_1/A dadda_fa_3_77_1/B dadda_fa_3_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_0/CIN dadda_fa_4_77_2/A sky130_fd_sc_hd__fa_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_54_0 dadda_fa_6_54_0/A dadda_fa_6_54_0/B dadda_fa_6_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_55_0/B dadda_fa_7_54_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater409 U$$622/A2 VGND VGND VPWR VPWR U$$574/A2 sky130_fd_sc_hd__buf_4
XFILLER_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4102 U$$4102/A U$$4109/A VGND VGND VPWR VPWR U$$4102/X sky130_fd_sc_hd__xor2_1
XFILLER_78_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4113 U$$4203/B U$$4113/B VGND VGND VPWR VPWR U$$4113/X sky130_fd_sc_hd__and2_1
XU$$4124 U$$4259/B1 U$$4140/A2 U$$4400/A1 U$$4140/B2 VGND VGND VPWR VPWR U$$4125/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4135 U$$4135/A U$$4215/B VGND VGND VPWR VPWR U$$4135/X sky130_fd_sc_hd__xor2_1
XU$$4146 U$$4418/B1 U$$4182/A2 U$$4285/A1 U$$4182/B2 VGND VGND VPWR VPWR U$$4147/A
+ sky130_fd_sc_hd__a22o_1
XU$$3401 U$$3401/A _665_/Q VGND VGND VPWR VPWR U$$3401/X sky130_fd_sc_hd__xor2_1
XFILLER_65_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4157 U$$4157/A U$$4183/B VGND VGND VPWR VPWR U$$4157/X sky130_fd_sc_hd__xor2_1
XU$$3412 U$$3412/A1 U$$3418/A2 U$$3412/B1 U$$3418/B2 VGND VGND VPWR VPWR U$$3413/A
+ sky130_fd_sc_hd__a22o_1
XU$$3423 U$$3423/A U$$3423/B VGND VGND VPWR VPWR U$$3423/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_113_2 dadda_fa_4_113_2/A dadda_fa_4_113_2/B dadda_fa_4_113_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_114_0/CIN dadda_fa_5_113_1/CIN sky130_fd_sc_hd__fa_1
XU$$4168 U$$4305/A1 U$$4226/A2 U$$4168/B1 U$$4226/B2 VGND VGND VPWR VPWR U$$4169/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3434 U$$3434/A U$$3478/B VGND VGND VPWR VPWR U$$3434/X sky130_fd_sc_hd__xor2_1
XU$$4179 U$$4179/A U$$4203/B VGND VGND VPWR VPWR U$$4179/X sky130_fd_sc_hd__xor2_1
XU$$2700 U$$2700/A U$$2708/B VGND VGND VPWR VPWR U$$2700/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3445 U$$3445/A1 U$$3479/A2 _559_/Q U$$3479/B2 VGND VGND VPWR VPWR U$$3446/A sky130_fd_sc_hd__a22o_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3456 U$$3456/A U$$3561/A VGND VGND VPWR VPWR U$$3456/X sky130_fd_sc_hd__xor2_1
XU$$2711 U$$2983/B1 U$$2607/X U$$2848/B1 U$$2608/X VGND VGND VPWR VPWR U$$2712/A sky130_fd_sc_hd__a22o_1
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2722 U$$2722/A U$$2730/B VGND VGND VPWR VPWR U$$2722/X sky130_fd_sc_hd__xor2_1
XFILLER_37_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3467 U$$4426/A1 U$$3545/A2 _570_/Q U$$3545/B2 VGND VGND VPWR VPWR U$$3468/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_106_1 dadda_fa_4_106_1/A dadda_fa_4_106_1/B dadda_fa_4_106_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/B dadda_fa_5_106_1/B sky130_fd_sc_hd__fa_1
XU$$2733 _613_/Q U$$2733/A2 _614_/Q U$$2733/B2 VGND VGND VPWR VPWR U$$2734/A sky130_fd_sc_hd__a22o_1
XFILLER_46_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3478 U$$3478/A U$$3478/B VGND VGND VPWR VPWR U$$3478/X sky130_fd_sc_hd__xor2_1
XU$$3489 _580_/Q U$$3519/A2 U$$4450/A1 U$$3519/B2 VGND VGND VPWR VPWR U$$3490/A sky130_fd_sc_hd__a22o_1
XU$$2744 U$$2742/Y _656_/Q _655_/Q U$$2743/X U$$2740/Y VGND VGND VPWR VPWR U$$2744/X
+ sky130_fd_sc_hd__a32o_4
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2755 U$$2755/A U$$2795/B VGND VGND VPWR VPWR U$$2755/X sky130_fd_sc_hd__xor2_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2766 U$$3312/B1 U$$2812/A2 U$$848/B1 U$$2812/B2 VGND VGND VPWR VPWR U$$2767/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2777 U$$2777/A U$$2827/B VGND VGND VPWR VPWR U$$2777/X sky130_fd_sc_hd__xor2_1
XFILLER_33_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2788 U$$596/A1 U$$2788/A2 U$$596/B1 U$$2788/B2 VGND VGND VPWR VPWR U$$2789/A sky130_fd_sc_hd__a22o_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2799 U$$2799/A U$$2839/B VGND VGND VPWR VPWR U$$2799/X sky130_fd_sc_hd__xor2_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_127_0 dadda_fa_7_127_0/A dadda_fa_7_127_0/B dadda_fa_7_127_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_127_0/COUT _423_/D sky130_fd_sc_hd__fa_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_72_0 dadda_fa_2_72_0/A dadda_fa_2_72_0/B dadda_fa_2_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_0/B dadda_fa_3_72_2/B sky130_fd_sc_hd__fa_1
XFILLER_29_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$706 final_adder.U$$706/A final_adder.U$$706/B VGND VGND VPWR VPWR
+ _252_/D sky130_fd_sc_hd__xor2_1
XFILLER_190_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater910 U$$4334/B VGND VGND VPWR VPWR U$$4322/B sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$717 final_adder.U$$717/A final_adder.U$$717/B VGND VGND VPWR VPWR
+ _263_/D sky130_fd_sc_hd__xor2_1
XFILLER_56_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater921 U$$4072/B VGND VGND VPWR VPWR U$$4044/B sky130_fd_sc_hd__buf_8
XFILLER_110_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$728 final_adder.U$$728/A final_adder.U$$728/B VGND VGND VPWR VPWR
+ _274_/D sky130_fd_sc_hd__xor2_4
Xrepeater932 U$$3933/B VGND VGND VPWR VPWR U$$3895/B sky130_fd_sc_hd__buf_8
Xfinal_adder.U$$739 final_adder.U$$739/A final_adder.U$$739/B VGND VGND VPWR VPWR
+ _285_/D sky130_fd_sc_hd__xor2_4
Xrepeater943 _671_/Q VGND VGND VPWR VPWR U$$3804/B sky130_fd_sc_hd__buf_6
Xrepeater954 U$$3663/B VGND VGND VPWR VPWR U$$3627/B sky130_fd_sc_hd__buf_8
XFILLER_56_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater965 _667_/Q VGND VGND VPWR VPWR U$$3562/A sky130_fd_sc_hd__buf_6
Xrepeater976 U$$3256/B VGND VGND VPWR VPWR U$$3218/B sky130_fd_sc_hd__buf_6
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater987 U$$3111/B VGND VGND VPWR VPWR U$$3077/B sky130_fd_sc_hd__buf_6
XFILLER_65_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater998 U$$3008/B VGND VGND VPWR VPWR U$$2982/B sky130_fd_sc_hd__buf_6
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3990 U$$3990/A U$$3994/B VGND VGND VPWR VPWR U$$3990/X sky130_fd_sc_hd__xor2_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_919 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_94_1 dadda_fa_4_94_1/A dadda_fa_4_94_1/B dadda_fa_4_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/B dadda_fa_5_94_1/B sky130_fd_sc_hd__fa_1
XFILLER_165_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_71_0 dadda_fa_7_71_0/A dadda_fa_7_71_0/B dadda_fa_7_71_0/CIN VGND VGND
+ VPWR VPWR _496_/D _367_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_87_0 dadda_fa_4_87_0/A dadda_fa_4_87_0/B dadda_fa_4_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/A dadda_fa_5_87_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_108_3 U$$4479/X input138/X dadda_fa_3_108_3/CIN VGND VGND VPWR VPWR dadda_fa_4_109_1/B
+ dadda_fa_4_108_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_161_640 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4391_1774 VGND VGND VPWR VPWR U$$4391_1774/HI U$$4391/B sky130_fd_sc_hd__conb_1
Xoutput270 _279_/Q VGND VGND VPWR VPWR o[111] sky130_fd_sc_hd__buf_2
XFILLER_0_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput281 _289_/Q VGND VGND VPWR VPWR o[121] sky130_fd_sc_hd__buf_2
Xoutput292 _184_/Q VGND VGND VPWR VPWR o[16] sky130_fd_sc_hd__buf_2
XFILLER_88_941 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4467_1812 VGND VGND VPWR VPWR U$$4467_1812/HI U$$4467/B sky130_fd_sc_hd__conb_1
XFILLER_130_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2007 U$$2007/A U$$2043/B VGND VGND VPWR VPWR U$$2007/X sky130_fd_sc_hd__xor2_1
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2018 U$$3386/B1 U$$2028/A2 U$$3388/B1 U$$2028/B2 VGND VGND VPWR VPWR U$$2019/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2029 U$$2029/A U$$2029/B VGND VGND VPWR VPWR U$$2029/X sky130_fd_sc_hd__xor2_1
XFILLER_210_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1306 U$$1306/A U$$1310/B VGND VGND VPWR VPWR U$$1306/X sky130_fd_sc_hd__xor2_1
XU$$1317 U$$3096/B1 U$$1355/A2 U$$2415/A1 U$$1355/B2 VGND VGND VPWR VPWR U$$1318/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1328 U$$1328/A U$$1332/B VGND VGND VPWR VPWR U$$1328/X sky130_fd_sc_hd__xor2_1
XU$$1339 U$$2435/A1 U$$1345/A2 U$$791/B1 U$$1345/B2 VGND VGND VPWR VPWR U$$1340/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_205_ _207_/CLK _205_/D VGND VGND VPWR VPWR _205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_51_5 dadda_fa_2_51_5/A dadda_fa_2_51_5/B dadda_fa_2_51_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_2/A dadda_fa_4_51_0/A sky130_fd_sc_hd__fa_1
XFILLER_93_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_955 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_44_4 dadda_fa_2_44_4/A dadda_fa_2_44_4/B dadda_fa_2_44_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_1/CIN dadda_fa_3_44_3/CIN sky130_fd_sc_hd__fa_1
XU$$3220 U$$3220/A U$$3256/B VGND VGND VPWR VPWR U$$3220/X sky130_fd_sc_hd__xor2_1
XFILLER_94_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_6_3_0 U$$13/X U$$146/X VGND VGND VPWR VPWR dadda_fa_7_4_0/B dadda_ha_6_3_0/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_24_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3231 U$$4464/A1 U$$3231/A2 U$$3779/B1 U$$3231/B2 VGND VGND VPWR VPWR U$$3232/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$13 _437_/Q _309_/Q VGND VGND VPWR VPWR final_adder.U$$141/B1 final_adder.U$$635/A
+ sky130_fd_sc_hd__ha_2
XU$$3242 U$$3242/A U$$3276/B VGND VGND VPWR VPWR U$$3242/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1050 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3253 U$$3388/B1 U$$3263/A2 U$$3253/B1 U$$3263/B2 VGND VGND VPWR VPWR U$$3254/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$24 _448_/Q _320_/Q VGND VGND VPWR VPWR final_adder.U$$519/B1 final_adder.U$$646/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$35 _459_/Q _331_/Q VGND VGND VPWR VPWR final_adder.U$$163/B1 final_adder.U$$657/A
+ sky130_fd_sc_hd__ha_1
XU$$3264 U$$3264/A U$$3272/B VGND VGND VPWR VPWR U$$3264/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_37_3 U$$1943/X U$$2076/X U$$2209/X VGND VGND VPWR VPWR dadda_fa_3_38_1/B
+ dadda_fa_3_37_3/B sky130_fd_sc_hd__fa_1
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$46 _470_/Q _342_/Q VGND VGND VPWR VPWR final_adder.U$$541/B1 final_adder.U$$668/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$57 _481_/Q _353_/Q VGND VGND VPWR VPWR final_adder.U$$185/B1 final_adder.U$$679/A
+ sky130_fd_sc_hd__ha_1
XU$$2530 U$$4035/B1 U$$2530/A2 U$$3902/A1 U$$2530/B2 VGND VGND VPWR VPWR U$$2531/A
+ sky130_fd_sc_hd__a22o_1
XU$$3275 U$$3412/A1 U$$3155/X U$$3412/B1 U$$3156/X VGND VGND VPWR VPWR U$$3276/A sky130_fd_sc_hd__a22o_1
XU$$3286 U$$3286/A U$$3286/B VGND VGND VPWR VPWR U$$3286/X sky130_fd_sc_hd__xor2_1
XFILLER_62_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2541 U$$2541/A U$$2541/B VGND VGND VPWR VPWR U$$2541/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2552 U$$908/A1 U$$2588/A2 U$$910/A1 U$$2588/B2 VGND VGND VPWR VPWR U$$2553/A sky130_fd_sc_hd__a22o_1
XU$$3297 U$$3297/A U$$3343/B VGND VGND VPWR VPWR U$$3297/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$68 _492_/Q _364_/Q VGND VGND VPWR VPWR final_adder.U$$563/B1 final_adder.U$$690/A
+ sky130_fd_sc_hd__ha_2
XFILLER_80_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$79 _503_/Q _375_/Q VGND VGND VPWR VPWR final_adder.U$$207/B1 final_adder.U$$701/A
+ sky130_fd_sc_hd__ha_1
XFILLER_181_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2563 U$$2563/A U$$2583/B VGND VGND VPWR VPWR U$$2563/X sky130_fd_sc_hd__xor2_1
XU$$2574 U$$4218/A1 U$$2580/A2 U$$4357/A1 U$$2580/B2 VGND VGND VPWR VPWR U$$2575/A
+ sky130_fd_sc_hd__a22o_1
XU$$1840 U$$1840/A U$$1844/B VGND VGND VPWR VPWR U$$1840/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2585 U$$2585/A U$$2603/A VGND VGND VPWR VPWR U$$2585/X sky130_fd_sc_hd__xor2_1
XU$$2596 _613_/Q U$$2600/A2 _614_/Q U$$2600/B2 VGND VGND VPWR VPWR U$$2597/A sky130_fd_sc_hd__a22o_1
XU$$1851 U$$3358/A1 U$$1851/A2 U$$2947/B1 U$$1851/B2 VGND VGND VPWR VPWR U$$1852/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1862 U$$1862/A U$$1870/B VGND VGND VPWR VPWR U$$1862/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1873 U$$3380/A1 U$$1907/A2 U$$2832/B1 U$$1907/B2 VGND VGND VPWR VPWR U$$1874/A
+ sky130_fd_sc_hd__a22o_1
XU$$1884 U$$1884/A U$$1884/B VGND VGND VPWR VPWR U$$1884/X sky130_fd_sc_hd__xor2_1
XU$$1895 U$$251/A1 U$$1915/A2 U$$251/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1896/A sky130_fd_sc_hd__a22o_1
XFILLER_148_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_868 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$503 final_adder.U$$8/SUM final_adder.U$$630/B final_adder.U$$8/COUT
+ VGND VGND VPWR VPWR final_adder.U$$631/B sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$525 final_adder.U$$652/A final_adder.U$$652/B final_adder.U$$525/B1
+ VGND VGND VPWR VPWR final_adder.U$$653/B sky130_fd_sc_hd__a21o_1
XFILLER_84_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater740 U$$3408/B2 VGND VGND VPWR VPWR U$$3404/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$547 final_adder.U$$674/A final_adder.U$$674/B final_adder.U$$547/B1
+ VGND VGND VPWR VPWR final_adder.U$$675/B sky130_fd_sc_hd__a21o_1
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater751 U$$3148/B2 VGND VGND VPWR VPWR U$$3066/B2 sky130_fd_sc_hd__buf_4
XFILLER_84_443 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater762 U$$3005/B2 VGND VGND VPWR VPWR U$$2959/B2 sky130_fd_sc_hd__buf_6
XFILLER_85_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$569 final_adder.U$$696/A final_adder.U$$696/B final_adder.U$$569/B1
+ VGND VGND VPWR VPWR final_adder.U$$697/B sky130_fd_sc_hd__a21o_1
XU$$408 U$$545/A1 U$$408/A2 U$$408/B1 U$$408/B2 VGND VGND VPWR VPWR U$$409/A sky130_fd_sc_hd__a22o_1
Xrepeater773 U$$408/B2 VGND VGND VPWR VPWR U$$392/B2 sky130_fd_sc_hd__buf_6
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$419 U$$828/B1 U$$447/A2 U$$556/B1 U$$447/B2 VGND VGND VPWR VPWR U$$420/A sky130_fd_sc_hd__a22o_1
Xrepeater784 U$$2663/B2 VGND VGND VPWR VPWR U$$2653/B2 sky130_fd_sc_hd__buf_4
Xrepeater795 U$$2471/X VGND VGND VPWR VPWR U$$2530/B2 sky130_fd_sc_hd__buf_4
XFILLER_198_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_47 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4497_1827 VGND VGND VPWR VPWR U$$4497_1827/HI U$$4497/B sky130_fd_sc_hd__conb_1
XFILLER_200_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1308 _601_/Q VGND VGND VPWR VPWR U$$3255/B1 sky130_fd_sc_hd__buf_4
XFILLER_154_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_113_1 U$$3824/X U$$3957/X U$$4090/X VGND VGND VPWR VPWR dadda_fa_4_114_2/A
+ dadda_fa_4_113_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater1319 U$$4214/A1 VGND VGND VPWR VPWR U$$4351/A1 sky130_fd_sc_hd__buf_4
XFILLER_114_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_106_0 U$$3544/X U$$3677/X U$$3810/X VGND VGND VPWR VPWR dadda_fa_4_107_0/B
+ dadda_fa_4_106_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_84_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_54_3 dadda_fa_3_54_3/A dadda_fa_3_54_3/B dadda_fa_3_54_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_1/B dadda_fa_4_54_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_125_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_47_2 dadda_fa_3_47_2/A dadda_fa_3_47_2/B dadda_fa_3_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_1/A dadda_fa_4_47_2/B sky130_fd_sc_hd__fa_1
XFILLER_208_438 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$920 U$$98/A1 U$$924/A2 U$$98/B1 U$$924/B2 VGND VGND VPWR VPWR U$$921/A sky130_fd_sc_hd__a22o_1
XU$$931 U$$931/A U$$935/B VGND VGND VPWR VPWR U$$931/X sky130_fd_sc_hd__xor2_1
XFILLER_18_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$942 U$$942/A1 U$$948/A2 U$$942/B1 U$$948/B2 VGND VGND VPWR VPWR U$$943/A sky130_fd_sc_hd__a22o_1
XU$$953 U$$953/A U$$958/A VGND VGND VPWR VPWR U$$953/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_17_0 dadda_fa_6_17_0/A dadda_fa_6_17_0/B dadda_fa_6_17_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_18_0/B dadda_fa_7_17_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_44_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$964 U$$962/B _629_/Q _630_/Q U$$959/Y VGND VGND VPWR VPWR U$$964/X sky130_fd_sc_hd__a22o_4
XU$$1103 U$$1103/A U$$1195/B VGND VGND VPWR VPWR U$$1103/X sky130_fd_sc_hd__xor2_1
XU$$1114 U$$18/A1 U$$1176/A2 U$$20/A1 U$$1176/B2 VGND VGND VPWR VPWR U$$1115/A sky130_fd_sc_hd__a22o_1
XU$$975 U$$16/A1 U$$979/A2 U$$18/A1 U$$979/B2 VGND VGND VPWR VPWR U$$976/A sky130_fd_sc_hd__a22o_1
XU$$1125 U$$1125/A U$$1151/B VGND VGND VPWR VPWR U$$1125/X sky130_fd_sc_hd__xor2_1
XU$$986 U$$986/A U$$998/B VGND VGND VPWR VPWR U$$986/X sky130_fd_sc_hd__xor2_1
XU$$1136 U$$2641/B1 U$$1146/A2 U$$2508/A1 U$$1146/B2 VGND VGND VPWR VPWR U$$1137/A
+ sky130_fd_sc_hd__a22o_1
XU$$997 U$$997/A1 U$$997/A2 U$$999/A1 U$$997/B2 VGND VGND VPWR VPWR U$$998/A sky130_fd_sc_hd__a22o_1
XFILLER_189_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1147 U$$1147/A U$$1147/B VGND VGND VPWR VPWR U$$1147/X sky130_fd_sc_hd__xor2_1
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_1018 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1158 U$$334/B1 U$$1190/A2 U$$201/A1 U$$1190/B2 VGND VGND VPWR VPWR U$$1159/A sky130_fd_sc_hd__a22o_1
XU$$1169 U$$1169/A U$$1177/B VGND VGND VPWR VPWR U$$1169/X sky130_fd_sc_hd__xor2_1
XFILLER_204_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_42_1 U$$2352/X U$$2485/X U$$2618/X VGND VGND VPWR VPWR dadda_fa_3_43_0/CIN
+ dadda_fa_3_42_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3050 U$$719/B1 U$$3054/A2 U$$3187/B1 U$$3054/B2 VGND VGND VPWR VPWR U$$3051/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_35_0 U$$343/X U$$476/X U$$609/X VGND VGND VPWR VPWR dadda_fa_3_36_0/B
+ dadda_fa_3_35_2/B sky130_fd_sc_hd__fa_1
XFILLER_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3061 U$$3061/A U$$3065/B VGND VGND VPWR VPWR U$$3061/X sky130_fd_sc_hd__xor2_1
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3072 U$$4305/A1 U$$3148/A2 U$$4168/B1 U$$3148/B2 VGND VGND VPWR VPWR U$$3073/A
+ sky130_fd_sc_hd__a22o_1
XU$$3083 U$$3083/A U$$3083/B VGND VGND VPWR VPWR U$$3083/X sky130_fd_sc_hd__xor2_1
XFILLER_179_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3094 U$$4053/A1 U$$3110/A2 U$$3096/A1 U$$3110/B2 VGND VGND VPWR VPWR U$$3095/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2360 U$$2360/A U$$2366/B VGND VGND VPWR VPWR U$$2360/X sky130_fd_sc_hd__xor2_1
XU$$2371 U$$2508/A1 U$$2423/A2 U$$2508/B1 U$$2423/B2 VGND VGND VPWR VPWR U$$2372/A
+ sky130_fd_sc_hd__a22o_1
XU$$2382 U$$2382/A U$$2388/B VGND VGND VPWR VPWR U$$2382/X sky130_fd_sc_hd__xor2_1
XU$$2393 U$$64/A1 U$$2395/A2 U$$66/A1 U$$2395/B2 VGND VGND VPWR VPWR U$$2394/A sky130_fd_sc_hd__a22o_1
XFILLER_34_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1670 U$$4410/A1 U$$1710/A2 U$$3042/A1 U$$1710/B2 VGND VGND VPWR VPWR U$$1671/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1681 U$$1681/A U$$1723/B VGND VGND VPWR VPWR U$$1681/X sky130_fd_sc_hd__xor2_1
XFILLER_179_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1692 U$$2786/B1 U$$1740/A2 U$$3475/A1 U$$1740/B2 VGND VGND VPWR VPWR U$$1693/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_87_3 U$$2841/X U$$2974/X U$$3107/X VGND VGND VPWR VPWR dadda_fa_2_88_4/A
+ dadda_fa_2_87_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_157_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_64_2 dadda_fa_4_64_2/A dadda_fa_4_64_2/B dadda_fa_4_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/CIN dadda_fa_5_64_1/CIN sky130_fd_sc_hd__fa_1
XTAP_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_57_1 dadda_fa_4_57_1/A dadda_fa_4_57_1/B dadda_fa_4_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/B dadda_fa_5_57_1/B sky130_fd_sc_hd__fa_1
XFILLER_170_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$300 final_adder.U$$300/A final_adder.U$$300/B VGND VGND VPWR VPWR
+ final_adder.U$$342/B sky130_fd_sc_hd__and2_2
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_34_0 dadda_fa_7_34_0/A dadda_fa_7_34_0/B dadda_fa_7_34_0/CIN VGND VGND
+ VPWR VPWR _459_/D _330_/D sky130_fd_sc_hd__fa_1
XFILLER_130_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$311 final_adder.U$$310/A final_adder.U$$237/X final_adder.U$$239/X
+ VGND VGND VPWR VPWR final_adder.U$$311/X sky130_fd_sc_hd__a21o_1
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$322 final_adder.U$$322/A final_adder.U$$322/B VGND VGND VPWR VPWR
+ final_adder.U$$322/X sky130_fd_sc_hd__and2_1
XFILLER_85_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$333 final_adder.U$$332/A final_adder.U$$281/X final_adder.U$$283/X
+ VGND VGND VPWR VPWR final_adder.U$$333/X sky130_fd_sc_hd__a21o_1
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$344 final_adder.U$$344/A final_adder.U$$344/B VGND VGND VPWR VPWR
+ final_adder.U$$364/B sky130_fd_sc_hd__and2_1
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$355 final_adder.U$$354/A final_adder.U$$325/X final_adder.U$$327/X
+ VGND VGND VPWR VPWR final_adder.U$$355/X sky130_fd_sc_hd__a21o_1
XU$$205 U$$614/B1 U$$217/A2 U$$344/A1 U$$217/B2 VGND VGND VPWR VPWR U$$206/A sky130_fd_sc_hd__a22o_1
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater570 U$$2145/A2 VGND VGND VPWR VPWR U$$2115/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$377 final_adder.U$$370/X final_adder.U$$654/B final_adder.U$$371/X
+ VGND VGND VPWR VPWR final_adder.U$$686/B sky130_fd_sc_hd__a21o_4
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater581 U$$2040/A2 VGND VGND VPWR VPWR U$$2052/A2 sky130_fd_sc_hd__buf_6
XFILLER_57_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$216 U$$216/A U$$216/B VGND VGND VPWR VPWR U$$216/X sky130_fd_sc_hd__xor2_1
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater592 U$$1648/X VGND VGND VPWR VPWR U$$1736/A2 sky130_fd_sc_hd__buf_4
XU$$227 U$$501/A1 U$$259/A2 U$$229/A1 U$$259/B2 VGND VGND VPWR VPWR U$$228/A sky130_fd_sc_hd__a22o_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$399 final_adder.U$$362/B final_adder.U$$702/B final_adder.U$$341/X
+ VGND VGND VPWR VPWR final_adder.U$$710/B sky130_fd_sc_hd__a21o_2
XU$$238 U$$238/A U$$250/B VGND VGND VPWR VPWR U$$238/X sky130_fd_sc_hd__xor2_1
XFILLER_55_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$249 U$$384/B1 U$$249/A2 U$$251/A1 U$$249/B2 VGND VGND VPWR VPWR U$$250/A sky130_fd_sc_hd__a22o_1
XFILLER_26_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_470_ _470_/CLK _470_/D VGND VGND VPWR VPWR _470_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1095 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1105 U$$1292/B VGND VGND VPWR VPWR U$$1296/B sky130_fd_sc_hd__buf_6
XFILLER_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1116 U$$1232/A VGND VGND VPWR VPWR U$$1225/B sky130_fd_sc_hd__buf_6
Xrepeater1127 U$$1078/B VGND VGND VPWR VPWR U$$1095/A sky130_fd_sc_hd__buf_8
Xrepeater1138 U$$796/B VGND VGND VPWR VPWR U$$726/B sky130_fd_sc_hd__buf_6
Xrepeater1149 U$$684/A VGND VGND VPWR VPWR U$$659/B sky130_fd_sc_hd__buf_6
XFILLER_5_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_75_1 U$$1221/X U$$1354/X U$$1487/X VGND VGND VPWR VPWR dadda_fa_1_76_8/B
+ dadda_fa_2_75_0/A sky130_fd_sc_hd__fa_1
XFILLER_49_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_52_0 dadda_fa_3_52_0/A dadda_fa_3_52_0/B dadda_fa_3_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_0/B dadda_fa_4_52_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_0_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_68_0 dadda_fa_0_68_0/A U$$409/X U$$542/X VGND VGND VPWR VPWR dadda_fa_1_69_5/CIN
+ dadda_fa_1_68_7/B sky130_fd_sc_hd__fa_1
XFILLER_208_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_668_ _674_/CLK _668_/D VGND VGND VPWR VPWR _668_/Q sky130_fd_sc_hd__dfxtp_1
XU$$750 U$$750/A U$$766/B VGND VGND VPWR VPWR U$$750/X sky130_fd_sc_hd__xor2_1
XU$$761 U$$896/B1 U$$765/A2 U$$761/B1 U$$765/B2 VGND VGND VPWR VPWR U$$762/A sky130_fd_sc_hd__a22o_1
XFILLER_95_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$772 U$$772/A U$$816/B VGND VGND VPWR VPWR U$$772/X sky130_fd_sc_hd__xor2_1
XFILLER_90_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$783 U$$98/A1 U$$783/A2 U$$98/B1 U$$783/B2 VGND VGND VPWR VPWR U$$784/A sky130_fd_sc_hd__a22o_1
XFILLER_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$794 U$$794/A U$$804/B VGND VGND VPWR VPWR U$$794/X sky130_fd_sc_hd__xor2_1
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_599_ _613_/CLK _599_/D VGND VGND VPWR VPWR _599_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_clk _369_/CLK VGND VGND VPWR VPWR _560_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_182_1176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_0 clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_2_97_2 U$$3127/X U$$3260/X U$$3393/X VGND VGND VPWR VPWR dadda_fa_3_98_1/A
+ dadda_fa_3_97_3/A sky130_fd_sc_hd__fa_1
XFILLER_67_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_74_1 dadda_fa_5_74_1/A dadda_fa_5_74_1/B dadda_fa_5_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_75_0/B dadda_fa_7_74_0/A sky130_fd_sc_hd__fa_1
XFILLER_67_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1650 _559_/Q VGND VGND VPWR VPWR U$$3310/A1 sky130_fd_sc_hd__buf_6
Xrepeater1661 U$$4404/A1 VGND VGND VPWR VPWR U$$4402/B1 sky130_fd_sc_hd__buf_6
Xrepeater1672 U$$3713/B1 VGND VGND VPWR VPWR U$$2345/A1 sky130_fd_sc_hd__buf_4
Xrepeater1683 U$$3163/B1 VGND VGND VPWR VPWR U$$562/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_5_67_0 dadda_fa_5_67_0/A dadda_fa_5_67_0/B dadda_fa_5_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_68_0/A dadda_fa_6_67_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1694 _554_/Q VGND VGND VPWR VPWR U$$3437/A1 sky130_fd_sc_hd__buf_4
XFILLER_28_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_66_8 dadda_fa_1_66_8/A dadda_fa_1_66_8/B dadda_fa_1_66_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_3/A dadda_fa_3_66_0/A sky130_fd_sc_hd__fa_2
XFILLER_6_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_59_7 dadda_fa_1_59_7/A dadda_fa_1_59_7/B dadda_fa_1_59_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_60_2/CIN dadda_fa_2_59_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_6_0 input223/X dadda_fa_6_6_0/B dadda_fa_6_6_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_7_7_0/B dadda_fa_7_6_0/CIN sky130_fd_sc_hd__fa_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2190 U$$2190/A U$$2191/A VGND VGND VPWR VPWR U$$2190/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_61_clk _535_/CLK VGND VGND VPWR VPWR _575_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_210_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_92_1 U$$2319/X U$$2452/X U$$2585/X VGND VGND VPWR VPWR dadda_fa_2_93_5/A
+ dadda_fa_2_92_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1069 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_85_0 U$$1506/Y U$$1640/X U$$1773/X VGND VGND VPWR VPWR dadda_fa_2_86_2/B
+ dadda_fa_2_85_4/B sky130_fd_sc_hd__fa_1
XFILLER_89_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4509 U$$4509/A U$$4509/B VGND VGND VPWR VPWR U$$4509/X sky130_fd_sc_hd__xor2_1
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$130 final_adder.U$$625/A final_adder.U$$624/A VGND VGND VPWR VPWR
+ final_adder.U$$130/X sky130_fd_sc_hd__and2_1
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3808 U$$3808/A U$$3836/A VGND VGND VPWR VPWR U$$3808/X sky130_fd_sc_hd__xor2_1
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3819 U$$4504/A1 U$$3703/X U$$4506/A1 U$$3704/X VGND VGND VPWR VPWR U$$3820/A sky130_fd_sc_hd__a22o_1
XFILLER_46_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$141 final_adder.U$$635/A final_adder.U$$507/B1 final_adder.U$$141/B1
+ VGND VGND VPWR VPWR final_adder.U$$141/X sky130_fd_sc_hd__a21o_1
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$152 final_adder.U$$647/A final_adder.U$$646/A VGND VGND VPWR VPWR
+ final_adder.U$$268/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$163 final_adder.U$$657/A final_adder.U$$529/B1 final_adder.U$$163/B1
+ VGND VGND VPWR VPWR final_adder.U$$163/X sky130_fd_sc_hd__a21o_1
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$174 final_adder.U$$669/A final_adder.U$$668/A VGND VGND VPWR VPWR
+ final_adder.U$$278/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$185 final_adder.U$$679/A final_adder.U$$551/B1 final_adder.U$$185/B1
+ VGND VGND VPWR VPWR final_adder.U$$185/X sky130_fd_sc_hd__a21o_1
XFILLER_205_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_522_ _523_/CLK _522_/D VGND VGND VPWR VPWR _522_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$196 final_adder.U$$691/A final_adder.U$$690/A VGND VGND VPWR VPWR
+ final_adder.U$$290/B sky130_fd_sc_hd__and2_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_5_126_0 dadda_ha_5_126_0/A U$$4382/X VGND VGND VPWR VPWR dadda_fa_7_127_0/A
+ dadda_fa_7_126_0/A sky130_fd_sc_hd__ha_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_453_ _469_/CLK _453_/D VGND VGND VPWR VPWR _453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_clk _535_/CLK VGND VGND VPWR VPWR _521_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_384_ _558_/CLK _384_/D VGND VGND VPWR VPWR _384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_303 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_84_0 dadda_fa_6_84_0/A dadda_fa_6_84_0/B dadda_fa_6_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_85_0/B dadda_fa_7_84_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput170 c[21] VGND VGND VPWR VPWR input170/X sky130_fd_sc_hd__clkbuf_4
Xinput181 c[31] VGND VGND VPWR VPWR input181/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput192 c[41] VGND VGND VPWR VPWR input192/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$580 U$$715/B1 U$$600/A2 U$$582/A1 U$$600/B2 VGND VGND VPWR VPWR U$$581/A sky130_fd_sc_hd__a22o_1
XFILLER_211_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$591 U$$591/A U$$669/B VGND VGND VPWR VPWR U$$591/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_43_clk _479_/CLK VGND VGND VPWR VPWR _503_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_177_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_98_0_1866 VGND VGND VPWR VPWR dadda_fa_2_98_0/A dadda_fa_2_98_0_1866/LO
+ sky130_fd_sc_hd__conb_1
Xrepeater1480 _580_/Q VGND VGND VPWR VPWR U$$4448/A1 sky130_fd_sc_hd__buf_8
XFILLER_99_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1491 _579_/Q VGND VGND VPWR VPWR U$$3624/A1 sky130_fd_sc_hd__buf_6
XFILLER_28_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_71_6 input225/X dadda_fa_1_71_6/B dadda_fa_1_71_6/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_72_2/B dadda_fa_2_71_5/B sky130_fd_sc_hd__fa_1
XFILLER_99_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_64_5 input217/X dadda_fa_1_64_5/B dadda_fa_1_64_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_65_2/A dadda_fa_2_64_5/A sky130_fd_sc_hd__fa_1
XFILLER_41_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_57_4 U$$2781/X U$$2914/X U$$3047/X VGND VGND VPWR VPWR dadda_fa_2_58_1/CIN
+ dadda_fa_2_57_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_27_2 dadda_fa_4_27_2/A dadda_fa_4_27_2/B dadda_fa_4_27_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/CIN dadda_fa_5_27_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_clk _479_/CLK VGND VGND VPWR VPWR _482_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_73 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4306 U$$4306/A U$$4348/B VGND VGND VPWR VPWR U$$4306/X sky130_fd_sc_hd__xor2_1
XU$$4317 _583_/Q U$$4327/A2 U$$4317/B1 U$$4319/B2 VGND VGND VPWR VPWR U$$4318/A sky130_fd_sc_hd__a22o_1
XFILLER_133_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4328 U$$4328/A U$$4334/B VGND VGND VPWR VPWR U$$4328/X sky130_fd_sc_hd__xor2_1
XFILLER_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4339 U$$4476/A1 U$$4251/X U$$4478/A1 U$$4345/B2 VGND VGND VPWR VPWR U$$4340/A
+ sky130_fd_sc_hd__a22o_1
XU$$3605 U$$3605/A U$$3609/B VGND VGND VPWR VPWR U$$3605/X sky130_fd_sc_hd__xor2_1
XU$$3616 U$$3753/A1 U$$3662/A2 U$$3618/A1 U$$3662/B2 VGND VGND VPWR VPWR U$$3617/A
+ sky130_fd_sc_hd__a22o_1
XU$$3627 U$$3627/A U$$3627/B VGND VGND VPWR VPWR U$$3627/X sky130_fd_sc_hd__xor2_1
XFILLER_46_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3638 U$$3638/A1 U$$3696/A2 U$$4462/A1 U$$3696/B2 VGND VGND VPWR VPWR U$$3639/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2904 U$$2904/A U$$2988/B VGND VGND VPWR VPWR U$$2904/X sky130_fd_sc_hd__xor2_1
XFILLER_93_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3649 U$$3649/A U$$3663/B VGND VGND VPWR VPWR U$$3649/X sky130_fd_sc_hd__xor2_1
XFILLER_34_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2915 U$$3187/B1 U$$2915/A2 U$$999/A1 U$$2915/B2 VGND VGND VPWR VPWR U$$2916/A
+ sky130_fd_sc_hd__a22o_1
XU$$2926 U$$2926/A U$$2928/B VGND VGND VPWR VPWR U$$2926/X sky130_fd_sc_hd__xor2_1
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_220 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2937 U$$4168/B1 U$$2973/A2 U$$4035/A1 U$$2973/B2 VGND VGND VPWR VPWR U$$2938/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_231 _188_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2948 U$$2948/A U$$2966/B VGND VGND VPWR VPWR U$$2948/X sky130_fd_sc_hd__xor2_1
XFILLER_93_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_505_ _507_/CLK _505_/D VGND VGND VPWR VPWR _505_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2959 U$$3916/B1 U$$2959/A2 U$$3783/A1 U$$2959/B2 VGND VGND VPWR VPWR U$$2960/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_980 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_22_1 U$$716/X U$$849/X U$$982/X VGND VGND VPWR VPWR dadda_fa_4_23_0/CIN
+ dadda_fa_4_22_2/A sky130_fd_sc_hd__fa_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_242 _192_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_253 _195_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_275 _212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clk _432_/CLK VGND VGND VPWR VPWR _463_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 _214_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_436_ _444_/CLK _436_/D VGND VGND VPWR VPWR _436_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_297 _233_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_367_ _496_/CLK _367_/D VGND VGND VPWR VPWR _367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_298_ _428_/CLK _298_/D VGND VGND VPWR VPWR _298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_81_5 dadda_fa_2_81_5/A dadda_fa_2_81_5/B dadda_fa_2_81_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_2/A dadda_fa_4_81_0/A sky130_fd_sc_hd__fa_2
XFILLER_181_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_74_4 dadda_fa_2_74_4/A dadda_fa_2_74_4/B dadda_fa_2_74_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/CIN dadda_fa_3_74_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_67_3 dadda_fa_2_67_3/A dadda_fa_2_67_3/B dadda_fa_2_67_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/B dadda_fa_3_67_3/B sky130_fd_sc_hd__fa_1
XFILLER_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_700 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_37_1 dadda_fa_5_37_1/A dadda_fa_5_37_1/B dadda_fa_5_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_38_0/B dadda_fa_7_37_0/A sky130_fd_sc_hd__fa_2
XFILLER_95_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk _432_/CLK VGND VGND VPWR VPWR _467_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_111_1 dadda_fa_5_111_1/A dadda_fa_5_111_1/B dadda_fa_5_111_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_112_0/B dadda_fa_7_111_0/A sky130_fd_sc_hd__fa_1
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_104_0 dadda_fa_5_104_0/A dadda_fa_5_104_0/B dadda_fa_5_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_105_0/A dadda_fa_6_104_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2198_1731 VGND VGND VPWR VPWR U$$2198_1731/HI U$$2198/A1 sky130_fd_sc_hd__conb_1
XFILLER_120_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_62_2 U$$3190/X U$$3323/X U$$3456/X VGND VGND VPWR VPWR dadda_fa_2_63_1/A
+ dadda_fa_2_62_4/A sky130_fd_sc_hd__fa_1
XFILLER_87_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_55_1 U$$1181/X U$$1314/X U$$1447/X VGND VGND VPWR VPWR dadda_fa_2_56_0/CIN
+ dadda_fa_2_55_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_41_1042 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_32_0 dadda_fa_4_32_0/A dadda_fa_4_32_0/B dadda_fa_4_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/A dadda_fa_5_32_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_48_0 U$$103/X U$$236/X U$$369/X VGND VGND VPWR VPWR dadda_fa_2_49_1/A
+ dadda_fa_2_48_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_500 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_221_ _482_/CLK _221_/D VGND VGND VPWR VPWR _221_/Q sky130_fd_sc_hd__dfxtp_1
Xdadda_fa_1_92_0_1860 VGND VGND VPWR VPWR dadda_fa_1_92_0/A dadda_fa_1_92_0_1860/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_211_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_502 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_84_3 dadda_fa_3_84_3/A dadda_fa_3_84_3/B dadda_fa_3_84_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_1/B dadda_fa_4_84_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_77_2 dadda_fa_3_77_2/A dadda_fa_3_77_2/B dadda_fa_3_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_1/A dadda_fa_4_77_2/B sky130_fd_sc_hd__fa_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_47_0 dadda_fa_6_47_0/A dadda_fa_6_47_0/B dadda_fa_6_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_48_0/B dadda_fa_7_47_0/CIN sky130_fd_sc_hd__fa_2
XU$$4103 U$$4238/B1 U$$4107/A2 U$$4105/A1 U$$4105/B2 VGND VGND VPWR VPWR U$$4104/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4114 U$$4112/Y _676_/Q _675_/Q U$$4113/X U$$4110/Y VGND VGND VPWR VPWR U$$4114/X
+ sky130_fd_sc_hd__a32o_4
XU$$4125 U$$4125/A U$$4141/B VGND VGND VPWR VPWR U$$4125/X sky130_fd_sc_hd__xor2_1
XFILLER_19_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4136 U$$4136/A1 U$$4140/A2 U$$4136/B1 U$$4140/B2 VGND VGND VPWR VPWR U$$4137/A
+ sky130_fd_sc_hd__a22o_1
XU$$4147 U$$4147/A U$$4183/B VGND VGND VPWR VPWR U$$4147/X sky130_fd_sc_hd__xor2_1
XU$$3402 U$$3539/A1 U$$3402/A2 _606_/Q U$$3402/B2 VGND VGND VPWR VPWR U$$3403/A sky130_fd_sc_hd__a22o_1
XU$$3413 U$$3413/A U$$3424/A VGND VGND VPWR VPWR U$$3413/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4158 U$$4158/A1 U$$4174/A2 U$$4160/A1 U$$4174/B2 VGND VGND VPWR VPWR U$$4159/A
+ sky130_fd_sc_hd__a22o_1
XU$$3424 U$$3424/A VGND VGND VPWR VPWR U$$3424/Y sky130_fd_sc_hd__inv_1
XU$$4169 U$$4169/A U$$4215/B VGND VGND VPWR VPWR U$$4169/X sky130_fd_sc_hd__xor2_1
XU$$3435 U$$3709/A1 U$$3479/A2 U$$3437/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3436/A
+ sky130_fd_sc_hd__a22o_1
XU$$2701 U$$4482/A1 U$$2607/X U$$4208/B1 U$$2608/X VGND VGND VPWR VPWR U$$2702/A sky130_fd_sc_hd__a22o_1
XU$$3446 U$$3446/A U$$3478/B VGND VGND VPWR VPWR U$$3446/X sky130_fd_sc_hd__xor2_1
XU$$3457 U$$4140/B1 U$$3559/A2 U$$4007/A1 U$$3559/B2 VGND VGND VPWR VPWR U$$3458/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2712 U$$2712/A U$$2739/A VGND VGND VPWR VPWR U$$2712/X sky130_fd_sc_hd__xor2_1
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2723 _608_/Q U$$2729/A2 U$$2725/A1 U$$2729/B2 VGND VGND VPWR VPWR U$$2724/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_106_2 dadda_fa_4_106_2/A dadda_fa_4_106_2/B dadda_fa_4_106_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/CIN dadda_fa_5_106_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3468 U$$3468/A U$$3506/B VGND VGND VPWR VPWR U$$3468/X sky130_fd_sc_hd__xor2_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3479 U$$4027/A1 U$$3479/A2 _576_/Q U$$3479/B2 VGND VGND VPWR VPWR U$$3480/A sky130_fd_sc_hd__a22o_1
XU$$2734 U$$2734/A U$$2734/B VGND VGND VPWR VPWR U$$2734/X sky130_fd_sc_hd__xor2_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2745 U$$2743/B _655_/Q _656_/Q U$$2740/Y VGND VGND VPWR VPWR U$$2745/X sky130_fd_sc_hd__a22o_4
XFILLER_61_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2756 U$$2756/A1 U$$2788/A2 U$$2756/B1 U$$2788/B2 VGND VGND VPWR VPWR U$$2757/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2767 U$$2767/A U$$2813/B VGND VGND VPWR VPWR U$$2767/X sky130_fd_sc_hd__xor2_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2778 U$$584/B1 U$$2812/A2 U$$4287/A1 U$$2812/B2 VGND VGND VPWR VPWR U$$2779/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2789 U$$2789/A U$$2795/B VGND VGND VPWR VPWR U$$2789/X sky130_fd_sc_hd__xor2_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_419_ _626_/CLK _419_/D VGND VGND VPWR VPWR _419_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1063 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_clk _442_/CLK VGND VGND VPWR VPWR _439_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_2_72_1 dadda_fa_2_72_1/A dadda_fa_2_72_1/B dadda_fa_2_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_0/CIN dadda_fa_3_72_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_110 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_644 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_65_0 dadda_fa_2_65_0/A dadda_fa_2_65_0/B dadda_fa_2_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_0/B dadda_fa_3_65_2/B sky130_fd_sc_hd__fa_1
Xrepeater900 U$$4496/B2 VGND VGND VPWR VPWR U$$4480/B2 sky130_fd_sc_hd__buf_6
XFILLER_64_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$707 final_adder.U$$707/A final_adder.U$$707/B VGND VGND VPWR VPWR
+ _253_/D sky130_fd_sc_hd__xor2_1
Xrepeater911 _679_/Q VGND VGND VPWR VPWR U$$4334/B sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$718 final_adder.U$$718/A final_adder.U$$718/B VGND VGND VPWR VPWR
+ _264_/D sky130_fd_sc_hd__xor2_1
XFILLER_29_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater922 U$$4036/B VGND VGND VPWR VPWR U$$3994/B sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$729 final_adder.U$$729/A final_adder.U$$729/B VGND VGND VPWR VPWR
+ _275_/D sky130_fd_sc_hd__xor2_4
XFILLER_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater933 U$$3943/B VGND VGND VPWR VPWR U$$3933/B sky130_fd_sc_hd__buf_6
XFILLER_99_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater944 U$$3816/B VGND VGND VPWR VPWR U$$3832/B sky130_fd_sc_hd__buf_6
Xrepeater955 U$$3671/B VGND VGND VPWR VPWR U$$3663/B sky130_fd_sc_hd__buf_8
Xrepeater966 _665_/Q VGND VGND VPWR VPWR U$$3397/B sky130_fd_sc_hd__buf_6
XFILLER_56_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater977 U$$3272/B VGND VGND VPWR VPWR U$$3256/B sky130_fd_sc_hd__buf_12
XFILLER_37_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater988 U$$3107/B VGND VGND VPWR VPWR U$$3111/B sky130_fd_sc_hd__buf_12
XFILLER_65_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater999 _659_/Q VGND VGND VPWR VPWR U$$3008/B sky130_fd_sc_hd__buf_6
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3980 U$$3980/A U$$4036/B VGND VGND VPWR VPWR U$$3980/X sky130_fd_sc_hd__xor2_1
XU$$3991 U$$4402/A1 U$$4005/A2 U$$4402/B1 U$$4005/B2 VGND VGND VPWR VPWR U$$3992/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_94_2 dadda_fa_4_94_2/A dadda_fa_4_94_2/B dadda_fa_4_94_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/CIN dadda_fa_5_94_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_180_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_87_1 dadda_fa_4_87_1/A dadda_fa_4_87_1/B dadda_fa_4_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/B dadda_fa_5_87_1/B sky130_fd_sc_hd__fa_1
XFILLER_133_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_64_0 dadda_fa_7_64_0/A dadda_fa_7_64_0/B dadda_fa_7_64_0/CIN VGND VGND
+ VPWR VPWR _489_/D _360_/D sky130_fd_sc_hd__fa_1
XFILLER_161_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput260 _270_/Q VGND VGND VPWR VPWR o[102] sky130_fd_sc_hd__buf_2
Xoutput271 _280_/Q VGND VGND VPWR VPWR o[112] sky130_fd_sc_hd__buf_2
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput282 _290_/Q VGND VGND VPWR VPWR o[122] sky130_fd_sc_hd__buf_2
Xoutput293 _185_/Q VGND VGND VPWR VPWR o[17] sky130_fd_sc_hd__buf_2
XFILLER_47_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_606 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2008 U$$2830/A1 U$$2038/A2 U$$3380/A1 U$$2038/B2 VGND VGND VPWR VPWR U$$2009/A
+ sky130_fd_sc_hd__a22o_1
XU$$2019 U$$2019/A U$$2029/B VGND VGND VPWR VPWR U$$2019/X sky130_fd_sc_hd__xor2_1
XFILLER_56_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1307 U$$74/A1 U$$1309/A2 U$$76/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1308/A sky130_fd_sc_hd__a22o_1
XFILLER_74_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1318 U$$1318/A U$$1356/B VGND VGND VPWR VPWR U$$1318/X sky130_fd_sc_hd__xor2_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1329 U$$2971/B1 U$$1237/X U$$2838/A1 U$$1238/X VGND VGND VPWR VPWR U$$1330/A sky130_fd_sc_hd__a22o_1
XFILLER_16_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_204_ _213_/CLK _204_/D VGND VGND VPWR VPWR _204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_82_0 dadda_fa_3_82_0/A dadda_fa_3_82_0/B dadda_fa_3_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_0/B dadda_fa_4_82_1/CIN sky130_fd_sc_hd__fa_1
XU$$4515_1836 VGND VGND VPWR VPWR U$$4515_1836/HI U$$4515/B sky130_fd_sc_hd__conb_1
XFILLER_48_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_387 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3210 U$$3210/A U$$3232/B VGND VGND VPWR VPWR U$$3210/X sky130_fd_sc_hd__xor2_1
XU$$3221 U$$3221/A1 U$$3263/A2 U$$3221/B1 U$$3263/B2 VGND VGND VPWR VPWR U$$3222/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_111_0 U$$4485/X input142/X dadda_fa_4_111_0/CIN VGND VGND VPWR VPWR dadda_fa_5_112_0/A
+ dadda_fa_5_111_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_44_5 dadda_fa_2_44_5/A dadda_fa_2_44_5/B dadda_fa_2_44_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_2/A dadda_fa_4_44_0/A sky130_fd_sc_hd__fa_1
XFILLER_19_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3232 U$$3232/A U$$3232/B VGND VGND VPWR VPWR U$$3232/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$14 _438_/Q _310_/Q VGND VGND VPWR VPWR final_adder.U$$509/B1 final_adder.U$$636/A
+ sky130_fd_sc_hd__ha_2
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$25 _449_/Q _321_/Q VGND VGND VPWR VPWR final_adder.U$$153/B1 final_adder.U$$647/A
+ sky130_fd_sc_hd__ha_2
XU$$3243 U$$3380/A1 U$$3283/A2 U$$4065/B1 U$$3283/B2 VGND VGND VPWR VPWR U$$3244/A
+ sky130_fd_sc_hd__a22o_1
XU$$3254 U$$3254/A U$$3256/B VGND VGND VPWR VPWR U$$3254/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$36 _460_/Q _332_/Q VGND VGND VPWR VPWR final_adder.U$$531/B1 final_adder.U$$658/A
+ sky130_fd_sc_hd__ha_1
XU$$3265 U$$3539/A1 U$$3273/A2 _606_/Q U$$3273/B2 VGND VGND VPWR VPWR U$$3266/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_37_4 U$$2342/X U$$2475/X input187/X VGND VGND VPWR VPWR dadda_fa_3_38_1/CIN
+ dadda_fa_3_37_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2520 U$$54/A1 U$$2524/A2 U$$56/A1 U$$2524/B2 VGND VGND VPWR VPWR U$$2521/A sky130_fd_sc_hd__a22o_1
XFILLER_98_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2531 U$$2531/A U$$2531/B VGND VGND VPWR VPWR U$$2531/X sky130_fd_sc_hd__xor2_1
XU$$3276 U$$3276/A U$$3276/B VGND VGND VPWR VPWR U$$3276/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$47 _471_/Q _343_/Q VGND VGND VPWR VPWR final_adder.U$$175/B1 final_adder.U$$669/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$58 _482_/Q _354_/Q VGND VGND VPWR VPWR final_adder.U$$553/B1 final_adder.U$$680/A
+ sky130_fd_sc_hd__ha_1
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2542 U$$3362/B1 U$$2566/A2 U$$3229/A1 U$$2566/B2 VGND VGND VPWR VPWR U$$2543/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_1095 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3287 U$$3288/A VGND VGND VPWR VPWR U$$3287/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$69 _493_/Q _365_/Q VGND VGND VPWR VPWR final_adder.U$$197/B1 final_adder.U$$691/A
+ sky130_fd_sc_hd__ha_2
XU$$2553 U$$2553/A U$$2597/B VGND VGND VPWR VPWR U$$2553/X sky130_fd_sc_hd__xor2_1
XU$$3298 U$$3709/A1 U$$3320/A2 U$$3437/A1 U$$3320/B2 VGND VGND VPWR VPWR U$$3299/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2564 U$$918/B1 U$$2566/A2 U$$3934/B1 U$$2566/B2 VGND VGND VPWR VPWR U$$2565/A
+ sky130_fd_sc_hd__a22o_1
XU$$2575 U$$2575/A U$$2583/B VGND VGND VPWR VPWR U$$2575/X sky130_fd_sc_hd__xor2_1
XU$$1830 U$$1830/A U$$1874/B VGND VGND VPWR VPWR U$$1830/X sky130_fd_sc_hd__xor2_1
XU$$1841 U$$3485/A1 U$$1843/A2 U$$1843/A1 U$$1843/B2 VGND VGND VPWR VPWR U$$1842/A
+ sky130_fd_sc_hd__a22o_1
XU$$2586 _608_/Q U$$2588/A2 U$$2586/B1 U$$2588/B2 VGND VGND VPWR VPWR U$$2587/A sky130_fd_sc_hd__a22o_1
XFILLER_22_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2597 U$$2597/A U$$2597/B VGND VGND VPWR VPWR U$$2597/X sky130_fd_sc_hd__xor2_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1852 U$$1852/A U$$1852/B VGND VGND VPWR VPWR U$$1852/X sky130_fd_sc_hd__xor2_1
XU$$1863 U$$3505/B1 U$$1785/X U$$358/A1 U$$1786/X VGND VGND VPWR VPWR U$$1864/A sky130_fd_sc_hd__a22o_1
XU$$1874 U$$1874/A U$$1874/B VGND VGND VPWR VPWR U$$1874/X sky130_fd_sc_hd__xor2_1
XU$$1885 U$$3253/B1 U$$1897/A2 U$$791/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1886/A
+ sky130_fd_sc_hd__a22o_1
XU$$1896 U$$1896/A U$$1917/A VGND VGND VPWR VPWR U$$1896/X sky130_fd_sc_hd__xor2_1
XFILLER_148_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_97_0 dadda_fa_5_97_0/A dadda_fa_5_97_0/B dadda_fa_5_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_98_0/A dadda_fa_6_97_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$515 final_adder.U$$642/A final_adder.U$$642/B final_adder.U$$515/B1
+ VGND VGND VPWR VPWR final_adder.U$$643/B sky130_fd_sc_hd__a21o_1
Xrepeater730 U$$3430/X VGND VGND VPWR VPWR U$$3537/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$537 final_adder.U$$664/A final_adder.U$$664/B final_adder.U$$537/B1
+ VGND VGND VPWR VPWR final_adder.U$$665/B sky130_fd_sc_hd__a21o_1
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater741 U$$3293/X VGND VGND VPWR VPWR U$$3408/B2 sky130_fd_sc_hd__buf_4
XFILLER_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater752 U$$3082/B2 VGND VGND VPWR VPWR U$$3046/B2 sky130_fd_sc_hd__buf_6
XFILLER_57_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater763 U$$3005/B2 VGND VGND VPWR VPWR U$$2997/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$559 final_adder.U$$686/A final_adder.U$$686/B final_adder.U$$559/B1
+ VGND VGND VPWR VPWR final_adder.U$$687/B sky130_fd_sc_hd__a21o_1
XFILLER_84_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater774 U$$279/X VGND VGND VPWR VPWR U$$408/B2 sky130_fd_sc_hd__clkbuf_8
XU$$409 U$$409/A U$$410/A VGND VGND VPWR VPWR U$$409/X sky130_fd_sc_hd__xor2_1
XFILLER_42_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater785 U$$2705/B2 VGND VGND VPWR VPWR U$$2663/B2 sky130_fd_sc_hd__buf_4
Xrepeater796 U$$2588/B2 VGND VGND VPWR VPWR U$$2600/B2 sky130_fd_sc_hd__buf_6
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_396 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1309 U$$3942/A1 VGND VGND VPWR VPWR U$$2435/A1 sky130_fd_sc_hd__buf_6
XFILLER_4_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_106_1 U$$3943/X U$$4076/X U$$4209/X VGND VGND VPWR VPWR dadda_fa_4_107_0/CIN
+ dadda_fa_4_106_2/A sky130_fd_sc_hd__fa_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_127_0 U$$4383/Y U$$4517/X input159/X VGND VGND VPWR VPWR dadda_fa_6_127_0/COUT
+ dadda_fa_7_127_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$271_1738 VGND VGND VPWR VPWR U$$271_1738/HI U$$271/B1 sky130_fd_sc_hd__conb_1
XFILLER_0_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_47_3 dadda_fa_3_47_3/A dadda_fa_3_47_3/B dadda_fa_3_47_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_1/B dadda_fa_4_47_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$910 U$$910/A1 U$$956/A2 U$$912/A1 U$$956/B2 VGND VGND VPWR VPWR U$$911/A sky130_fd_sc_hd__a22o_1
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$921 U$$921/A U$$925/B VGND VGND VPWR VPWR U$$921/X sky130_fd_sc_hd__xor2_1
XFILLER_29_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$932 U$$932/A1 U$$826/X U$$934/A1 U$$827/X VGND VGND VPWR VPWR U$$933/A sky130_fd_sc_hd__a22o_1
XFILLER_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$943 U$$943/A U$$951/B VGND VGND VPWR VPWR U$$943/X sky130_fd_sc_hd__xor2_1
XU$$954 U$$954/A1 U$$956/A2 U$$956/A1 U$$956/B2 VGND VGND VPWR VPWR U$$955/A sky130_fd_sc_hd__a22o_1
XFILLER_16_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$965 U$$965/A1 U$$995/A2 U$$967/A1 U$$995/B2 VGND VGND VPWR VPWR U$$966/A sky130_fd_sc_hd__a22o_1
XU$$1104 U$$967/A1 U$$1194/A2 U$$969/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1105/A sky130_fd_sc_hd__a22o_1
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$976 U$$976/A U$$980/B VGND VGND VPWR VPWR U$$976/X sky130_fd_sc_hd__xor2_1
XU$$1115 U$$1115/A U$$1177/B VGND VGND VPWR VPWR U$$1115/X sky130_fd_sc_hd__xor2_1
XFILLER_203_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1126 U$$989/A1 U$$1194/A2 U$$991/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1127/A sky130_fd_sc_hd__a22o_1
XU$$987 U$$987/A1 U$$997/A2 U$$30/A1 U$$997/B2 VGND VGND VPWR VPWR U$$988/A sky130_fd_sc_hd__a22o_1
XFILLER_204_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1137 U$$1137/A U$$1147/B VGND VGND VPWR VPWR U$$1137/X sky130_fd_sc_hd__xor2_1
XU$$998 U$$998/A U$$998/B VGND VGND VPWR VPWR U$$998/X sky130_fd_sc_hd__xor2_1
XFILLER_204_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1148 U$$52/A1 U$$1176/A2 U$$52/B1 U$$1176/B2 VGND VGND VPWR VPWR U$$1149/A sky130_fd_sc_hd__a22o_1
XFILLER_188_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1159 U$$1159/A U$$1191/B VGND VGND VPWR VPWR U$$1159/X sky130_fd_sc_hd__xor2_1
XFILLER_31_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_42_2 U$$2751/X U$$2884/X U$$2928/B VGND VGND VPWR VPWR dadda_fa_3_43_1/A
+ dadda_fa_3_42_3/A sky130_fd_sc_hd__fa_1
XFILLER_66_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3040 U$$4410/A1 U$$3082/A2 U$$3042/A1 U$$3082/B2 VGND VGND VPWR VPWR U$$3041/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_371 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3051 U$$3051/A U$$3077/B VGND VGND VPWR VPWR U$$3051/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_1 U$$742/X U$$875/X U$$1008/X VGND VGND VPWR VPWR dadda_fa_3_36_0/CIN
+ dadda_fa_3_35_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3062 U$$4432/A1 U$$3066/A2 U$$4434/A1 U$$3066/B2 VGND VGND VPWR VPWR U$$3063/A
+ sky130_fd_sc_hd__a22o_1
XU$$3073 U$$3073/A U$$3107/B VGND VGND VPWR VPWR U$$3073/X sky130_fd_sc_hd__xor2_1
XU$$3084 U$$3221/A1 U$$3110/A2 U$$3221/B1 U$$3110/B2 VGND VGND VPWR VPWR U$$3085/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_330 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_12_0 input160/X dadda_fa_5_12_0/B dadda_fa_5_12_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_6_13_0/A dadda_fa_6_12_0/CIN sky130_fd_sc_hd__fa_1
XU$$3095 U$$3095/A U$$3111/B VGND VGND VPWR VPWR U$$3095/X sky130_fd_sc_hd__xor2_1
XFILLER_35_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2350 U$$2350/A U$$2400/B VGND VGND VPWR VPWR U$$2350/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_28_0 U$$63/X U$$196/X U$$329/X VGND VGND VPWR VPWR dadda_fa_3_29_1/CIN
+ dadda_fa_3_28_3/A sky130_fd_sc_hd__fa_1
XFILLER_35_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2361 U$$3181/B1 U$$2367/A2 U$$3046/B1 U$$2367/B2 VGND VGND VPWR VPWR U$$2362/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2372 U$$2372/A U$$2418/B VGND VGND VPWR VPWR U$$2372/X sky130_fd_sc_hd__xor2_1
XFILLER_35_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2383 U$$3342/A1 U$$2387/A2 U$$4027/B1 U$$2387/B2 VGND VGND VPWR VPWR U$$2384/A
+ sky130_fd_sc_hd__a22o_1
XU$$2394 U$$2394/A U$$2400/B VGND VGND VPWR VPWR U$$2394/X sky130_fd_sc_hd__xor2_1
XFILLER_201_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1660 U$$2756/A1 U$$1736/A2 U$$2756/B1 U$$1736/B2 VGND VGND VPWR VPWR U$$1661/A
+ sky130_fd_sc_hd__a22o_1
XU$$1671 U$$1671/A U$$1711/B VGND VGND VPWR VPWR U$$1671/X sky130_fd_sc_hd__xor2_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1682 U$$997/A1 U$$1740/A2 U$$999/A1 U$$1740/B2 VGND VGND VPWR VPWR U$$1683/A sky130_fd_sc_hd__a22o_1
XFILLER_210_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1693 U$$1693/A U$$1723/B VGND VGND VPWR VPWR U$$1693/X sky130_fd_sc_hd__xor2_1
XFILLER_194_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_87_4 U$$3240/X U$$3373/X U$$3506/X VGND VGND VPWR VPWR dadda_fa_2_88_4/B
+ dadda_fa_3_87_0/A sky130_fd_sc_hd__fa_1
XFILLER_118_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_57_2 dadda_fa_4_57_2/A dadda_fa_4_57_2/B dadda_fa_4_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/CIN dadda_fa_5_57_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$301 final_adder.U$$300/A final_adder.U$$217/X final_adder.U$$219/X
+ VGND VGND VPWR VPWR final_adder.U$$301/X sky130_fd_sc_hd__a21o_2
XFILLER_170_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$312 final_adder.U$$312/A final_adder.U$$312/B VGND VGND VPWR VPWR
+ final_adder.U$$348/B sky130_fd_sc_hd__and2_1
XFILLER_40_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$323 final_adder.U$$322/A final_adder.U$$261/X final_adder.U$$263/X
+ VGND VGND VPWR VPWR final_adder.U$$323/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$334 final_adder.U$$334/A final_adder.U$$334/B VGND VGND VPWR VPWR
+ final_adder.U$$358/A sky130_fd_sc_hd__and2_1
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$345 final_adder.U$$344/A final_adder.U$$305/X final_adder.U$$307/X
+ VGND VGND VPWR VPWR final_adder.U$$345/X sky130_fd_sc_hd__a21o_1
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$356 final_adder.U$$356/A final_adder.U$$356/B VGND VGND VPWR VPWR
+ final_adder.U$$370/B sky130_fd_sc_hd__and2_1
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater560 U$$2248/A2 VGND VGND VPWR VPWR U$$2242/A2 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_7_27_0 dadda_fa_7_27_0/A dadda_fa_7_27_0/B dadda_fa_7_27_0/CIN VGND VGND
+ VPWR VPWR _452_/D _323_/D sky130_fd_sc_hd__fa_1
XU$$206 U$$206/A U$$216/B VGND VGND VPWR VPWR U$$206/X sky130_fd_sc_hd__xor2_1
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater571 U$$2169/A2 VGND VGND VPWR VPWR U$$2145/A2 sky130_fd_sc_hd__buf_6
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater582 U$$1922/X VGND VGND VPWR VPWR U$$2040/A2 sky130_fd_sc_hd__buf_8
XU$$217 U$$900/B1 U$$217/A2 U$$82/A1 U$$217/B2 VGND VGND VPWR VPWR U$$218/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$389 final_adder.U$$364/X final_adder.U$$718/B final_adder.U$$365/X
+ VGND VGND VPWR VPWR final_adder.U$$734/B sky130_fd_sc_hd__a21o_4
Xrepeater593 U$$1718/A2 VGND VGND VPWR VPWR U$$1710/A2 sky130_fd_sc_hd__buf_6
XU$$228 U$$228/A U$$232/B VGND VGND VPWR VPWR U$$228/X sky130_fd_sc_hd__xor2_1
XFILLER_57_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$239 U$$648/B1 U$$249/A2 U$$650/B1 U$$249/B2 VGND VGND VPWR VPWR U$$240/A sky130_fd_sc_hd__a22o_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1069 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_79 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1106 U$$1288/B VGND VGND VPWR VPWR U$$1292/B sky130_fd_sc_hd__buf_6
Xrepeater1117 U$$1209/B VGND VGND VPWR VPWR U$$1232/A sky130_fd_sc_hd__buf_12
Xrepeater1128 _631_/Q VGND VGND VPWR VPWR U$$1078/B sky130_fd_sc_hd__buf_6
XFILLER_49_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1139 U$$804/B VGND VGND VPWR VPWR U$$760/B sky130_fd_sc_hd__buf_8
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_52_1 dadda_fa_3_52_1/A dadda_fa_3_52_1/B dadda_fa_3_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_0/CIN dadda_fa_4_52_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_0_68_1 U$$675/X U$$808/X U$$941/X VGND VGND VPWR VPWR dadda_fa_1_69_6/A
+ dadda_fa_1_68_7/CIN sky130_fd_sc_hd__fa_1
XTAP_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_45_0 dadda_fa_3_45_0/A dadda_fa_3_45_0/B dadda_fa_3_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_0/B dadda_fa_4_45_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$740 U$$740/A U$$748/B VGND VGND VPWR VPWR U$$740/X sky130_fd_sc_hd__xor2_1
XFILLER_1_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$751 U$$66/A1 U$$759/A2 U$$66/B1 U$$759/B2 VGND VGND VPWR VPWR U$$752/A sky130_fd_sc_hd__a22o_1
X_667_ _674_/CLK _667_/D VGND VGND VPWR VPWR _667_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_205_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$762 U$$762/A U$$766/B VGND VGND VPWR VPWR U$$762/X sky130_fd_sc_hd__xor2_1
XU$$773 U$$910/A1 U$$783/A2 U$$912/A1 U$$783/B2 VGND VGND VPWR VPWR U$$774/A sky130_fd_sc_hd__a22o_1
XU$$784 U$$784/A U$$816/B VGND VGND VPWR VPWR U$$784/X sky130_fd_sc_hd__xor2_1
XFILLER_56_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$795 U$$932/A1 U$$795/A2 U$$934/A1 U$$795/B2 VGND VGND VPWR VPWR U$$796/A sky130_fd_sc_hd__a22o_1
X_598_ _598_/CLK _598_/D VGND VGND VPWR VPWR _598_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_147_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_2_98_5 U$$4326/X U$$4459/X VGND VGND VPWR VPWR dadda_fa_3_99_2/B dadda_fa_4_98_0/A
+ sky130_fd_sc_hd__ha_1
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_102_0 dadda_fa_7_102_0/A dadda_fa_7_102_0/B dadda_fa_7_102_0/CIN VGND
+ VGND VPWR VPWR _527_/D _398_/D sky130_fd_sc_hd__fa_1
XFILLER_32_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 _566_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_2_97_3 U$$3526/X U$$3659/X U$$3792/X VGND VGND VPWR VPWR dadda_fa_3_98_1/B
+ dadda_fa_3_97_3/B sky130_fd_sc_hd__fa_1
XFILLER_160_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1640 U$$3584/B1 VGND VGND VPWR VPWR U$$435/A1 sky130_fd_sc_hd__buf_4
XFILLER_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1651 _559_/Q VGND VGND VPWR VPWR U$$2625/A1 sky130_fd_sc_hd__buf_6
Xrepeater1662 _558_/Q VGND VGND VPWR VPWR U$$4404/A1 sky130_fd_sc_hd__buf_6
XFILLER_153_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1673 U$$3713/B1 VGND VGND VPWR VPWR U$$973/B1 sky130_fd_sc_hd__buf_4
XFILLER_141_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1684 U$$4259/B1 VGND VGND VPWR VPWR U$$3163/B1 sky130_fd_sc_hd__buf_8
XFILLER_193_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_67_1 dadda_fa_5_67_1/A dadda_fa_5_67_1/B dadda_fa_5_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_68_0/B dadda_fa_7_67_0/A sky130_fd_sc_hd__fa_1
XFILLER_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1695 U$$2611/B1 VGND VGND VPWR VPWR U$$8/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_59_8 dadda_fa_1_59_8/A dadda_fa_1_59_8/B dadda_fa_1_59_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_60_3/A dadda_fa_3_59_0/A sky130_fd_sc_hd__fa_2
XFILLER_27_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_106_0 dadda_fa_2_106_0/A U$$3012/X U$$3145/X VGND VGND VPWR VPWR dadda_fa_3_107_3/B
+ dadda_fa_3_106_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_81_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2180 U$$2180/A U$$2186/B VGND VGND VPWR VPWR U$$2180/X sky130_fd_sc_hd__xor2_1
XU$$2191 U$$2191/A VGND VGND VPWR VPWR U$$2191/Y sky130_fd_sc_hd__inv_1
XFILLER_34_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1490 U$$2721/B1 U$$1500/A2 U$$2725/A1 U$$1500/B2 VGND VGND VPWR VPWR U$$1491/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_438 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_780 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_85_1 U$$1906/X U$$2039/X U$$2172/X VGND VGND VPWR VPWR dadda_fa_2_86_2/CIN
+ dadda_fa_2_85_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_116_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_62_0 dadda_fa_4_62_0/A dadda_fa_4_62_0/B dadda_fa_4_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/A dadda_fa_5_62_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_78_0 U$$1227/X U$$1360/X U$$1493/X VGND VGND VPWR VPWR dadda_fa_2_79_0/B
+ dadda_fa_2_78_3/B sky130_fd_sc_hd__fa_1
XFILLER_132_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_731 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$120 _544_/Q _416_/Q VGND VGND VPWR VPWR final_adder.U$$615/B1 final_adder.U$$742/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$131 final_adder.U$$625/A final_adder.U$$497/B1 final_adder.U$$3/COUT
+ VGND VGND VPWR VPWR final_adder.U$$131/X sky130_fd_sc_hd__a21o_1
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3809 U$$4355/B1 U$$3823/A2 U$$4222/A1 U$$3823/B2 VGND VGND VPWR VPWR U$$3810/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$142 final_adder.U$$637/A final_adder.U$$636/A VGND VGND VPWR VPWR
+ final_adder.U$$262/A sky130_fd_sc_hd__and2_1
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$153 final_adder.U$$647/A final_adder.U$$519/B1 final_adder.U$$153/B1
+ VGND VGND VPWR VPWR final_adder.U$$153/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$164 final_adder.U$$659/A final_adder.U$$658/A VGND VGND VPWR VPWR
+ final_adder.U$$274/B sky130_fd_sc_hd__and2_1
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$175 final_adder.U$$669/A final_adder.U$$541/B1 final_adder.U$$175/B1
+ VGND VGND VPWR VPWR final_adder.U$$175/X sky130_fd_sc_hd__a21o_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$186 final_adder.U$$681/A final_adder.U$$680/A VGND VGND VPWR VPWR
+ final_adder.U$$284/A sky130_fd_sc_hd__and2_1
Xrepeater390 U$$1093/A2 VGND VGND VPWR VPWR U$$1089/A2 sky130_fd_sc_hd__buf_4
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_521_ _521_/CLK _521_/D VGND VGND VPWR VPWR _521_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$197 final_adder.U$$691/A final_adder.U$$563/B1 final_adder.U$$197/B1
+ VGND VGND VPWR VPWR final_adder.U$$197/X sky130_fd_sc_hd__a21o_1
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_452_ _469_/CLK _452_/D VGND VGND VPWR VPWR _452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_383_ _572_/CLK _383_/D VGND VGND VPWR VPWR _383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_77_0 dadda_fa_6_77_0/A dadda_fa_6_77_0/B dadda_fa_6_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_78_0/B dadda_fa_7_77_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput160 c[12] VGND VGND VPWR VPWR input160/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput171 c[22] VGND VGND VPWR VPWR input171/X sky130_fd_sc_hd__buf_2
XFILLER_209_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput182 c[32] VGND VGND VPWR VPWR input182/X sky130_fd_sc_hd__buf_2
XFILLER_37_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput193 c[42] VGND VGND VPWR VPWR input193/X sky130_fd_sc_hd__clkbuf_1
XTAP_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$570 U$$707/A1 U$$574/A2 U$$22/B1 U$$574/B2 VGND VGND VPWR VPWR U$$571/A sky130_fd_sc_hd__a22o_1
XFILLER_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$581 U$$581/A U$$613/B VGND VGND VPWR VPWR U$$581/X sky130_fd_sc_hd__xor2_1
XFILLER_63_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$592 U$$42/B1 U$$622/A2 U$$729/B1 U$$622/B2 VGND VGND VPWR VPWR U$$593/A sky130_fd_sc_hd__a22o_1
XFILLER_32_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_95_0 U$$2591/X U$$2724/X U$$2857/X VGND VGND VPWR VPWR dadda_fa_3_96_0/B
+ dadda_fa_3_95_2/B sky130_fd_sc_hd__fa_1
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1470 U$$4450/A1 VGND VGND VPWR VPWR U$$3626/B1 sky130_fd_sc_hd__buf_6
Xrepeater1481 U$$4446/B1 VGND VGND VPWR VPWR U$$4035/B1 sky130_fd_sc_hd__buf_4
XFILLER_99_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1492 U$$745/A1 VGND VGND VPWR VPWR U$$882/A1 sky130_fd_sc_hd__buf_6
XFILLER_141_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_71_7 dadda_fa_1_71_7/A dadda_fa_1_71_7/B dadda_fa_1_71_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_72_2/CIN dadda_fa_2_71_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_64_6 dadda_fa_1_64_6/A dadda_fa_1_64_6/B dadda_fa_1_64_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_2/B dadda_fa_2_64_5/B sky130_fd_sc_hd__fa_1
XFILLER_74_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_57_5 U$$3180/X U$$3313/X U$$3446/X VGND VGND VPWR VPWR dadda_fa_2_58_2/A
+ dadda_fa_2_57_5/A sky130_fd_sc_hd__fa_1
XFILLER_41_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_94_0 dadda_fa_7_94_0/A dadda_fa_7_94_0/B dadda_fa_7_94_0/CIN VGND VGND
+ VPWR VPWR _519_/D _390_/D sky130_fd_sc_hd__fa_2
XFILLER_195_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1055 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4307 U$$4444/A1 U$$4251/X U$$4444/B1 U$$4345/B2 VGND VGND VPWR VPWR U$$4308/A
+ sky130_fd_sc_hd__a22o_1
XU$$4318 U$$4318/A U$$4322/B VGND VGND VPWR VPWR U$$4318/X sky130_fd_sc_hd__xor2_1
XU$$4329 U$$4466/A1 U$$4335/A2 U$$4468/A1 U$$4333/B2 VGND VGND VPWR VPWR U$$4330/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3606 U$$4291/A1 U$$3628/A2 U$$4293/A1 U$$3628/B2 VGND VGND VPWR VPWR U$$3607/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3617 U$$3617/A U$$3627/B VGND VGND VPWR VPWR U$$3617/X sky130_fd_sc_hd__xor2_1
XFILLER_92_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3628 U$$4176/A1 U$$3628/A2 U$$4176/B1 U$$3628/B2 VGND VGND VPWR VPWR U$$3629/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3639 U$$3639/A _669_/Q VGND VGND VPWR VPWR U$$3639/X sky130_fd_sc_hd__xor2_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2905 U$$3042/A1 U$$2959/A2 U$$3042/B1 U$$2959/B2 VGND VGND VPWR VPWR U$$2906/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2916 U$$2916/A U$$2916/B VGND VGND VPWR VPWR U$$2916/X sky130_fd_sc_hd__xor2_1
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2927 U$$4434/A1 U$$2929/A2 U$$4436/A1 U$$2929/B2 VGND VGND VPWR VPWR U$$2928/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2938 U$$2938/A U$$2972/B VGND VGND VPWR VPWR U$$2938/X sky130_fd_sc_hd__xor2_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 _188_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_504_ _504_/CLK _504_/D VGND VGND VPWR VPWR _504_/Q sky130_fd_sc_hd__dfxtp_1
XU$$2949 U$$3221/B1 U$$2959/A2 U$$3088/A1 U$$2959/B2 VGND VGND VPWR VPWR U$$2950/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_22_2 U$$1115/X U$$1248/X U$$1381/X VGND VGND VPWR VPWR dadda_fa_4_23_1/A
+ dadda_fa_4_22_2/B sky130_fd_sc_hd__fa_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_243 _193_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_254 _195_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 _212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_287 _214_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_435_ _435_/CLK _435_/D VGND VGND VPWR VPWR _435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_298 _233_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_444 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_366_ _495_/CLK _366_/D VGND VGND VPWR VPWR _366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_297_ _431_/CLK _297_/D VGND VGND VPWR VPWR _297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_74_5 dadda_fa_2_74_5/A dadda_fa_2_74_5/B dadda_fa_2_74_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_2/A dadda_fa_4_74_0/A sky130_fd_sc_hd__fa_1
XFILLER_96_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_271 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_67_4 dadda_fa_2_67_4/A dadda_fa_2_67_4/B dadda_fa_2_67_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/CIN dadda_fa_3_67_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_104_1 dadda_fa_5_104_1/A dadda_fa_5_104_1/B dadda_fa_5_104_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_105_0/B dadda_fa_7_104_0/A sky130_fd_sc_hd__fa_1
XFILLER_172_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_62_3 U$$3589/X U$$3722/X U$$3855/X VGND VGND VPWR VPWR dadda_fa_2_63_1/B
+ dadda_fa_2_62_4/B sky130_fd_sc_hd__fa_1
XFILLER_59_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_55_2 U$$1580/X U$$1713/X U$$1846/X VGND VGND VPWR VPWR dadda_fa_2_56_1/A
+ dadda_fa_2_55_4/A sky130_fd_sc_hd__fa_1
XFILLER_132_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_32_1 dadda_fa_4_32_1/A dadda_fa_4_32_1/B dadda_fa_4_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/B dadda_fa_5_32_1/B sky130_fd_sc_hd__fa_1
XFILLER_103_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_48_1 U$$502/X U$$635/X U$$768/X VGND VGND VPWR VPWR dadda_fa_2_49_1/B
+ dadda_fa_2_48_4/A sky130_fd_sc_hd__fa_1
XFILLER_27_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_25_0 dadda_fa_4_25_0/A dadda_fa_4_25_0/B dadda_fa_4_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/A dadda_fa_5_25_1/A sky130_fd_sc_hd__fa_1
XFILLER_103_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_220_ _482_/CLK _220_/D VGND VGND VPWR VPWR _220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_978 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_77_3 dadda_fa_3_77_3/A dadda_fa_3_77_3/B dadda_fa_3_77_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_1/B dadda_fa_4_77_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4104 U$$4104/A U$$4109/A VGND VGND VPWR VPWR U$$4104/X sky130_fd_sc_hd__xor2_1
XFILLER_24_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4115 U$$4113/B _675_/Q _676_/Q U$$4110/Y VGND VGND VPWR VPWR U$$4115/X sky130_fd_sc_hd__a22o_2
XU$$4126 U$$4400/A1 U$$4140/A2 U$$4402/A1 U$$4140/B2 VGND VGND VPWR VPWR U$$4127/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4137 U$$4137/A U$$4141/B VGND VGND VPWR VPWR U$$4137/X sky130_fd_sc_hd__xor2_1
XU$$4148 U$$4285/A1 U$$4182/A2 U$$4287/A1 U$$4182/B2 VGND VGND VPWR VPWR U$$4149/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_14_0 U$$35/X U$$168/X VGND VGND VPWR VPWR dadda_fa_4_15_2/B dadda_ha_3_14_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$3403 U$$3403/A _665_/Q VGND VGND VPWR VPWR U$$3403/X sky130_fd_sc_hd__xor2_1
XU$$4159 U$$4159/A U$$4175/B VGND VGND VPWR VPWR U$$4159/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3414 U$$4510/A1 U$$3292/X U$$3551/B1 U$$3293/X VGND VGND VPWR VPWR U$$3415/A sky130_fd_sc_hd__a22o_1
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3425 U$$3425/A VGND VGND VPWR VPWR U$$3425/Y sky130_fd_sc_hd__inv_1
XFILLER_19_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3436 U$$3436/A U$$3490/B VGND VGND VPWR VPWR U$$3436/X sky130_fd_sc_hd__xor2_1
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2702 U$$2702/A U$$2739/A VGND VGND VPWR VPWR U$$2702/X sky130_fd_sc_hd__xor2_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3447 _559_/Q U$$3497/A2 U$$3447/B1 U$$3497/B2 VGND VGND VPWR VPWR U$$3448/A sky130_fd_sc_hd__a22o_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2713 _603_/Q U$$2733/A2 U$$3674/A1 U$$2733/B2 VGND VGND VPWR VPWR U$$2714/A sky130_fd_sc_hd__a22o_1
XU$$3458 U$$3458/A U$$3561/A VGND VGND VPWR VPWR U$$3458/X sky130_fd_sc_hd__xor2_1
XU$$2724 U$$2724/A U$$2730/B VGND VGND VPWR VPWR U$$2724/X sky130_fd_sc_hd__xor2_1
XU$$3469 _570_/Q U$$3545/A2 U$$4430/A1 U$$3545/B2 VGND VGND VPWR VPWR U$$3470/A sky130_fd_sc_hd__a22o_1
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2735 U$$3283/A1 U$$2607/X U$$2872/B1 U$$2608/X VGND VGND VPWR VPWR U$$2736/A sky130_fd_sc_hd__a22o_1
XFILLER_34_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2746 U$$2746/A1 U$$2788/A2 U$$2746/B1 U$$2788/B2 VGND VGND VPWR VPWR U$$2747/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2757 U$$2757/A U$$2795/B VGND VGND VPWR VPWR U$$2757/X sky130_fd_sc_hd__xor2_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2768 U$$3042/A1 U$$2814/A2 U$$3042/B1 U$$2814/B2 VGND VGND VPWR VPWR U$$2769/A
+ sky130_fd_sc_hd__a22o_1
XU$$2779 U$$2779/A U$$2827/B VGND VGND VPWR VPWR U$$2779/X sky130_fd_sc_hd__xor2_1
XFILLER_61_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_418_ _547_/CLK _418_/D VGND VGND VPWR VPWR _418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_349_ _476_/CLK _349_/D VGND VGND VPWR VPWR _349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_72_2 dadda_fa_2_72_2/A dadda_fa_2_72_2/B dadda_fa_2_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/A dadda_fa_3_72_3/A sky130_fd_sc_hd__fa_1
XFILLER_68_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_65_1 dadda_fa_2_65_1/A dadda_fa_2_65_1/B dadda_fa_2_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_0/CIN dadda_fa_3_65_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater901 U$$4389/X VGND VGND VPWR VPWR U$$4516/B2 sky130_fd_sc_hd__clkbuf_4
Xfinal_adder.U$$708 final_adder.U$$708/A final_adder.U$$708/B VGND VGND VPWR VPWR
+ _254_/D sky130_fd_sc_hd__xor2_1
Xrepeater912 U$$4197/B VGND VGND VPWR VPWR U$$4183/B sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$719 final_adder.U$$719/A final_adder.U$$719/B VGND VGND VPWR VPWR
+ _265_/D sky130_fd_sc_hd__xor2_1
Xrepeater923 U$$4096/B VGND VGND VPWR VPWR U$$4036/B sky130_fd_sc_hd__buf_6
Xdadda_fa_5_42_0 dadda_fa_5_42_0/A dadda_fa_5_42_0/B dadda_fa_5_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_43_0/A dadda_fa_6_42_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater934 U$$3949/B VGND VGND VPWR VPWR U$$3965/B sky130_fd_sc_hd__buf_12
Xdadda_fa_2_58_0 dadda_fa_2_58_0/A dadda_fa_2_58_0/B dadda_fa_2_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_0/B dadda_fa_3_58_2/B sky130_fd_sc_hd__fa_1
Xrepeater945 U$$3836/A VGND VGND VPWR VPWR U$$3816/B sky130_fd_sc_hd__buf_6
XFILLER_204_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater956 _669_/Q VGND VGND VPWR VPWR U$$3671/B sky130_fd_sc_hd__buf_12
Xrepeater967 U$$3363/B VGND VGND VPWR VPWR U$$3357/B sky130_fd_sc_hd__buf_12
XFILLER_83_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater978 U$$3276/B VGND VGND VPWR VPWR U$$3272/B sky130_fd_sc_hd__buf_6
Xrepeater989 U$$3145/B VGND VGND VPWR VPWR U$$3107/B sky130_fd_sc_hd__buf_6
XFILLER_204_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3970 U$$4105/B1 U$$3970/A2 U$$3970/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3971/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3981 U$$4392/A1 U$$4005/A2 U$$4394/A1 U$$4005/B2 VGND VGND VPWR VPWR U$$3982/A
+ sky130_fd_sc_hd__a22o_1
XU$$3992 U$$3992/A U$$3994/B VGND VGND VPWR VPWR U$$3992/X sky130_fd_sc_hd__xor2_1
XFILLER_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4425_1791 VGND VGND VPWR VPWR U$$4425_1791/HI U$$4425/B sky130_fd_sc_hd__conb_1
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_87_2 dadda_fa_4_87_2/A dadda_fa_4_87_2/B dadda_fa_4_87_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/CIN dadda_fa_5_87_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput261 _271_/Q VGND VGND VPWR VPWR o[103] sky130_fd_sc_hd__buf_2
Xdadda_fa_7_57_0 dadda_fa_7_57_0/A dadda_fa_7_57_0/B dadda_fa_7_57_0/CIN VGND VGND
+ VPWR VPWR _482_/D _353_/D sky130_fd_sc_hd__fa_1
XFILLER_121_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput272 _281_/Q VGND VGND VPWR VPWR o[113] sky130_fd_sc_hd__buf_2
XFILLER_88_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput283 _291_/Q VGND VGND VPWR VPWR o[123] sky130_fd_sc_hd__buf_2
Xoutput294 _186_/Q VGND VGND VPWR VPWR o[18] sky130_fd_sc_hd__buf_2
XFILLER_58_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_47 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3148_1746 VGND VGND VPWR VPWR U$$3148_1746/HI U$$3148/B1 sky130_fd_sc_hd__conb_1
Xdadda_fa_1_60_0 U$$1989/X U$$2122/X U$$2255/X VGND VGND VPWR VPWR dadda_fa_2_61_0/B
+ dadda_fa_2_60_3/B sky130_fd_sc_hd__fa_1
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2009 U$$2009/A U$$2011/B VGND VGND VPWR VPWR U$$2009/X sky130_fd_sc_hd__xor2_1
XFILLER_90_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1308 U$$1308/A U$$1310/B VGND VGND VPWR VPWR U$$1308/X sky130_fd_sc_hd__xor2_1
XFILLER_167_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1319 U$$2415/A1 U$$1355/A2 U$$634/B1 U$$1355/B2 VGND VGND VPWR VPWR U$$1320/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_203_ _213_/CLK _203_/D VGND VGND VPWR VPWR _203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_82_1 dadda_fa_3_82_1/A dadda_fa_3_82_1/B dadda_fa_3_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_0/CIN dadda_fa_4_82_2/A sky130_fd_sc_hd__fa_1
XFILLER_180_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_75_0 dadda_fa_3_75_0/A dadda_fa_3_75_0/B dadda_fa_3_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_0/B dadda_fa_4_75_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_139_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3200 U$$3200/A U$$3236/B VGND VGND VPWR VPWR U$$3200/X sky130_fd_sc_hd__xor2_1
XU$$3211 _578_/Q U$$3231/A2 U$$3896/B1 U$$3231/B2 VGND VGND VPWR VPWR U$$3212/A sky130_fd_sc_hd__a22o_1
XFILLER_19_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3222 U$$3222/A U$$3256/B VGND VGND VPWR VPWR U$$3222/X sky130_fd_sc_hd__xor2_1
XFILLER_171_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_111_1 dadda_fa_4_111_1/A dadda_fa_4_111_1/B dadda_fa_4_111_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_112_0/B dadda_fa_5_111_1/B sky130_fd_sc_hd__fa_1
XFILLER_93_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3233 U$$3779/B1 U$$3283/A2 U$$3646/A1 U$$3283/B2 VGND VGND VPWR VPWR U$$3234/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$15 _439_/Q _311_/Q VGND VGND VPWR VPWR final_adder.U$$143/B1 final_adder.U$$637/A
+ sky130_fd_sc_hd__ha_2
XU$$3244 U$$3244/A U$$3276/B VGND VGND VPWR VPWR U$$3244/X sky130_fd_sc_hd__xor2_1
XU$$3255 _600_/Q U$$3263/A2 U$$3255/B1 U$$3263/B2 VGND VGND VPWR VPWR U$$3256/A sky130_fd_sc_hd__a22o_1
XU$$2510 U$$4154/A1 U$$2550/A2 U$$4154/B1 U$$2550/B2 VGND VGND VPWR VPWR U$$2511/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$26 _450_/Q _322_/Q VGND VGND VPWR VPWR final_adder.U$$521/B1 final_adder.U$$648/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$37 _461_/Q _333_/Q VGND VGND VPWR VPWR final_adder.U$$165/B1 final_adder.U$$659/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_2_37_5 dadda_fa_2_37_5/A dadda_fa_2_37_5/B dadda_fa_2_37_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_38_2/A dadda_fa_4_37_0/A sky130_fd_sc_hd__fa_2
XFILLER_4_1187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_104_0 dadda_fa_4_104_0/A dadda_fa_4_104_0/B dadda_fa_4_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/A dadda_fa_5_104_1/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$48 _472_/Q _344_/Q VGND VGND VPWR VPWR final_adder.U$$543/B1 final_adder.U$$670/A
+ sky130_fd_sc_hd__ha_1
XFILLER_185_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3266 U$$3266/A U$$3272/B VGND VGND VPWR VPWR U$$3266/X sky130_fd_sc_hd__xor2_1
XFILLER_19_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2521 U$$2521/A U$$2541/B VGND VGND VPWR VPWR U$$2521/X sky130_fd_sc_hd__xor2_1
XFILLER_206_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2532 U$$3902/A1 U$$2470/X U$$3902/B1 U$$2471/X VGND VGND VPWR VPWR U$$2533/A sky130_fd_sc_hd__a22o_1
XU$$3277 U$$3412/B1 U$$3283/A2 U$$3551/B1 U$$3283/B2 VGND VGND VPWR VPWR U$$3278/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$59 _483_/Q _355_/Q VGND VGND VPWR VPWR final_adder.U$$187/B1 final_adder.U$$681/A
+ sky130_fd_sc_hd__ha_1
XU$$3288 U$$3288/A VGND VGND VPWR VPWR U$$3288/Y sky130_fd_sc_hd__inv_1
XU$$2543 U$$2543/A U$$2567/B VGND VGND VPWR VPWR U$$2543/X sky130_fd_sc_hd__xor2_1
XU$$2554 U$$4061/A1 U$$2588/A2 U$$3652/A1 U$$2588/B2 VGND VGND VPWR VPWR U$$2555/A
+ sky130_fd_sc_hd__a22o_1
XU$$3299 U$$3299/A U$$3363/B VGND VGND VPWR VPWR U$$3299/X sky130_fd_sc_hd__xor2_1
XFILLER_179_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1820 U$$1820/A U$$1820/B VGND VGND VPWR VPWR U$$1820/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2565 U$$2565/A U$$2567/B VGND VGND VPWR VPWR U$$2565/X sky130_fd_sc_hd__xor2_1
XU$$1831 U$$50/A1 U$$1851/A2 U$$52/A1 U$$1851/B2 VGND VGND VPWR VPWR U$$1832/A sky130_fd_sc_hd__a22o_1
XFILLER_62_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2576 U$$3807/B1 U$$2580/A2 U$$3674/A1 U$$2580/B2 VGND VGND VPWR VPWR U$$2577/A
+ sky130_fd_sc_hd__a22o_1
XU$$1842 U$$1842/A U$$1844/B VGND VGND VPWR VPWR U$$1842/X sky130_fd_sc_hd__xor2_1
XU$$2587 U$$2587/A U$$2597/B VGND VGND VPWR VPWR U$$2587/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2598 _614_/Q U$$2600/A2 U$$2872/B1 U$$2600/B2 VGND VGND VPWR VPWR U$$2599/A sky130_fd_sc_hd__a22o_1
XFILLER_61_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1853 U$$2947/B1 U$$1907/A2 U$$896/A1 U$$1907/B2 VGND VGND VPWR VPWR U$$1854/A
+ sky130_fd_sc_hd__a22o_1
XU$$1864 U$$1864/A U$$1870/B VGND VGND VPWR VPWR U$$1864/X sky130_fd_sc_hd__xor2_1
XU$$1875 U$$2832/B1 U$$1909/A2 U$$3245/B1 U$$1909/B2 VGND VGND VPWR VPWR U$$1876/A
+ sky130_fd_sc_hd__a22o_1
XU$$1886 U$$1886/A U$$1917/A VGND VGND VPWR VPWR U$$1886/X sky130_fd_sc_hd__xor2_1
XFILLER_148_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1897 U$$2171/A1 U$$1897/A2 U$$392/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1898/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_97_1 dadda_fa_5_97_1/A dadda_fa_5_97_1/B dadda_fa_5_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_98_0/B dadda_fa_7_97_0/A sky130_fd_sc_hd__fa_1
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$505 final_adder.U$$632/A final_adder.U$$632/B final_adder.U$$505/B1
+ VGND VGND VPWR VPWR final_adder.U$$633/B sky130_fd_sc_hd__a21o_1
XFILLER_111_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater720 U$$3696/B2 VGND VGND VPWR VPWR U$$3636/B2 sky130_fd_sc_hd__buf_8
Xfinal_adder.U$$527 final_adder.U$$654/A final_adder.U$$654/B final_adder.U$$527/B1
+ VGND VGND VPWR VPWR final_adder.U$$655/B sky130_fd_sc_hd__a21o_1
Xrepeater731 U$$3545/B2 VGND VGND VPWR VPWR U$$3559/B2 sky130_fd_sc_hd__buf_4
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater742 U$$3285/B2 VGND VGND VPWR VPWR U$$3209/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_111_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$549 final_adder.U$$676/A final_adder.U$$676/B final_adder.U$$549/B1
+ VGND VGND VPWR VPWR final_adder.U$$677/B sky130_fd_sc_hd__a21o_1
Xrepeater753 U$$3110/B2 VGND VGND VPWR VPWR U$$3082/B2 sky130_fd_sc_hd__buf_8
Xrepeater764 U$$3005/B2 VGND VGND VPWR VPWR U$$2981/B2 sky130_fd_sc_hd__buf_12
XFILLER_84_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater775 U$$2812/B2 VGND VGND VPWR VPWR U$$2814/B2 sky130_fd_sc_hd__buf_6
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater786 U$$2707/B2 VGND VGND VPWR VPWR U$$2705/B2 sky130_fd_sc_hd__buf_6
Xrepeater797 U$$2580/B2 VGND VGND VPWR VPWR U$$2588/B2 sky130_fd_sc_hd__buf_6
XFILLER_37_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4490 U$$928/A1 U$$4388/X U$$4490/B1 U$$4496/B2 VGND VGND VPWR VPWR U$$4491/A sky130_fd_sc_hd__a22o_1
XFILLER_53_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2052_1728 VGND VGND VPWR VPWR U$$2052_1728/HI U$$2052/B1 sky130_fd_sc_hd__conb_1
XFILLER_80_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_92_0 dadda_fa_4_92_0/A dadda_fa_4_92_0/B dadda_fa_4_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/A dadda_fa_5_92_1/A sky130_fd_sc_hd__fa_1
XFILLER_14_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_106_2 U$$4342/X U$$4475/X input136/X VGND VGND VPWR VPWR dadda_fa_4_107_1/A
+ dadda_fa_4_106_2/B sky130_fd_sc_hd__fa_1
XFILLER_106_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_892 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$900 U$$900/A1 U$$906/A2 U$$900/B1 U$$906/B2 VGND VGND VPWR VPWR U$$901/A sky130_fd_sc_hd__a22o_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$911 U$$911/A U$$958/A VGND VGND VPWR VPWR U$$911/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_80_0_1854 VGND VGND VPWR VPWR dadda_fa_1_80_0/A dadda_fa_1_80_0_1854/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_63_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$922 U$$922/A1 U$$924/A2 U$$924/A1 U$$924/B2 VGND VGND VPWR VPWR U$$923/A sky130_fd_sc_hd__a22o_1
XU$$933 U$$933/A U$$935/B VGND VGND VPWR VPWR U$$933/X sky130_fd_sc_hd__xor2_1
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$944 U$$944/A1 U$$948/A2 U$$944/B1 U$$948/B2 VGND VGND VPWR VPWR U$$945/A sky130_fd_sc_hd__a22o_1
XU$$955 U$$955/A U$$958/A VGND VGND VPWR VPWR U$$955/X sky130_fd_sc_hd__xor2_1
XFILLER_204_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1105 U$$1105/A U$$1195/B VGND VGND VPWR VPWR U$$1105/X sky130_fd_sc_hd__xor2_1
XU$$966 U$$966/A U$$994/B VGND VGND VPWR VPWR U$$966/X sky130_fd_sc_hd__xor2_1
XU$$977 U$$18/A1 U$$979/A2 U$$20/A1 U$$979/B2 VGND VGND VPWR VPWR U$$978/A sky130_fd_sc_hd__a22o_1
XFILLER_44_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1116 U$$429/B1 U$$1150/A2 U$$22/A1 U$$1150/B2 VGND VGND VPWR VPWR U$$1117/A sky130_fd_sc_hd__a22o_1
XU$$1127 U$$1127/A U$$1195/B VGND VGND VPWR VPWR U$$1127/X sky130_fd_sc_hd__xor2_1
XU$$988 U$$988/A U$$998/B VGND VGND VPWR VPWR U$$988/X sky130_fd_sc_hd__xor2_1
XU$$1138 U$$2508/A1 U$$1146/A2 U$$2508/B1 U$$1146/B2 VGND VGND VPWR VPWR U$$1139/A
+ sky130_fd_sc_hd__a22o_1
XU$$999 U$$999/A1 U$$999/A2 U$$999/B1 U$$999/B2 VGND VGND VPWR VPWR U$$999/X sky130_fd_sc_hd__a22o_1
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1149 U$$1149/A U$$1177/B VGND VGND VPWR VPWR U$$1149/X sky130_fd_sc_hd__xor2_1
XFILLER_188_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_29_3 U$$1262/X U$$1395/X VGND VGND VPWR VPWR dadda_fa_3_30_2/B dadda_fa_4_29_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_42_3 input193/X dadda_fa_2_42_3/B dadda_fa_2_42_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_43_1/B dadda_fa_3_42_3/B sky130_fd_sc_hd__fa_1
XU$$3030 U$$3578/A1 U$$3046/A2 U$$3578/B1 U$$3046/B2 VGND VGND VPWR VPWR U$$3031/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3041 U$$3041/A U$$3083/B VGND VGND VPWR VPWR U$$3041/X sky130_fd_sc_hd__xor2_1
XFILLER_82_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3052 U$$3187/B1 U$$3054/A2 U$$3054/A1 U$$3054/B2 VGND VGND VPWR VPWR U$$3053/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_35_2 U$$1141/X U$$1274/X U$$1407/X VGND VGND VPWR VPWR dadda_fa_3_36_1/A
+ dadda_fa_3_35_3/A sky130_fd_sc_hd__fa_1
XFILLER_19_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3063 U$$3063/A U$$3065/B VGND VGND VPWR VPWR U$$3063/X sky130_fd_sc_hd__xor2_1
XU$$3074 U$$4031/B1 U$$3082/A2 U$$3896/B1 U$$3082/B2 VGND VGND VPWR VPWR U$$3075/A
+ sky130_fd_sc_hd__a22o_1
XU$$2340 U$$2340/A U$$2418/B VGND VGND VPWR VPWR U$$2340/X sky130_fd_sc_hd__xor2_1
XU$$3085 U$$3085/A U$$3111/B VGND VGND VPWR VPWR U$$3085/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_12_1 dadda_fa_5_12_1/A dadda_fa_5_12_1/B dadda_ha_4_12_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_13_0/B dadda_fa_7_12_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_28_1 U$$462/X U$$595/X U$$728/X VGND VGND VPWR VPWR dadda_fa_3_29_2/A
+ dadda_fa_3_28_3/B sky130_fd_sc_hd__fa_1
XFILLER_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2351 U$$2625/A1 U$$2395/A2 U$$435/A1 U$$2395/B2 VGND VGND VPWR VPWR U$$2352/A
+ sky130_fd_sc_hd__a22o_1
XU$$3096 U$$3096/A1 U$$3110/A2 U$$3096/B1 U$$3110/B2 VGND VGND VPWR VPWR U$$3097/A
+ sky130_fd_sc_hd__a22o_1
XU$$2362 U$$2362/A U$$2366/B VGND VGND VPWR VPWR U$$2362/X sky130_fd_sc_hd__xor2_1
XU$$2373 U$$2508/B1 U$$2423/A2 U$$2375/A1 U$$2423/B2 VGND VGND VPWR VPWR U$$2374/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2384 U$$2384/A U$$2388/B VGND VGND VPWR VPWR U$$2384/X sky130_fd_sc_hd__xor2_1
XU$$1650 U$$1650/A1 U$$1684/A2 U$$2746/B1 U$$1684/B2 VGND VGND VPWR VPWR U$$1651/A
+ sky130_fd_sc_hd__a22o_1
XU$$2395 U$$66/A1 U$$2395/A2 U$$66/B1 U$$2395/B2 VGND VGND VPWR VPWR U$$2396/A sky130_fd_sc_hd__a22o_1
XU$$1661 U$$1661/A U$$1687/B VGND VGND VPWR VPWR U$$1661/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1672 U$$3042/A1 U$$1710/A2 U$$3042/B1 U$$1710/B2 VGND VGND VPWR VPWR U$$1673/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1683 U$$1683/A U$$1723/B VGND VGND VPWR VPWR U$$1683/X sky130_fd_sc_hd__xor2_1
XU$$1694 U$$3475/A1 U$$1740/A2 U$$3475/B1 U$$1740/B2 VGND VGND VPWR VPWR U$$1695/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$302 final_adder.U$$302/A final_adder.U$$302/B VGND VGND VPWR VPWR
+ final_adder.U$$342/A sky130_fd_sc_hd__and2_1
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$313 final_adder.U$$312/A final_adder.U$$241/X final_adder.U$$243/X
+ VGND VGND VPWR VPWR final_adder.U$$313/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$324 final_adder.U$$324/A final_adder.U$$324/B VGND VGND VPWR VPWR
+ final_adder.U$$354/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$335 final_adder.U$$334/A final_adder.U$$285/X final_adder.U$$287/X
+ VGND VGND VPWR VPWR final_adder.U$$335/X sky130_fd_sc_hd__a21o_1
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$346 final_adder.U$$346/A final_adder.U$$346/B VGND VGND VPWR VPWR
+ final_adder.U$$364/A sky130_fd_sc_hd__and2_2
Xrepeater550 U$$2470/X VGND VGND VPWR VPWR U$$2580/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$357 final_adder.U$$356/A final_adder.U$$329/X final_adder.U$$331/X
+ VGND VGND VPWR VPWR final_adder.U$$357/X sky130_fd_sc_hd__a21o_1
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater561 U$$2302/A2 VGND VGND VPWR VPWR U$$2248/A2 sky130_fd_sc_hd__buf_6
XU$$207 U$$344/A1 U$$217/A2 U$$72/A1 U$$217/B2 VGND VGND VPWR VPWR U$$208/A sky130_fd_sc_hd__a22o_1
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater572 U$$2059/X VGND VGND VPWR VPWR U$$2169/A2 sky130_fd_sc_hd__buf_4
Xrepeater583 U$$1785/X VGND VGND VPWR VPWR U$$1859/A2 sky130_fd_sc_hd__buf_6
XFILLER_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$218 U$$218/A U$$232/B VGND VGND VPWR VPWR U$$218/X sky130_fd_sc_hd__xor2_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$229 U$$229/A1 U$$259/A2 U$$94/A1 U$$259/B2 VGND VGND VPWR VPWR U$$230/A sky130_fd_sc_hd__a22o_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater594 U$$1768/A2 VGND VGND VPWR VPWR U$$1718/A2 sky130_fd_sc_hd__buf_4
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1001 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1107 U$$1332/B VGND VGND VPWR VPWR U$$1288/B sky130_fd_sc_hd__buf_6
XFILLER_14_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_111_0 U$$3287/Y U$$3421/X U$$3554/X VGND VGND VPWR VPWR dadda_fa_4_112_1/A
+ dadda_fa_4_111_2/A sky130_fd_sc_hd__fa_1
Xrepeater1118 U$$1203/B VGND VGND VPWR VPWR U$$1209/B sky130_fd_sc_hd__buf_6
Xrepeater1129 U$$929/B VGND VGND VPWR VPWR U$$859/B sky130_fd_sc_hd__clkbuf_8
XFILLER_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_52_2 dadda_fa_3_52_2/A dadda_fa_3_52_2/B dadda_fa_3_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_1/A dadda_fa_4_52_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_0_68_2 U$$1074/X U$$1207/X U$$1340/X VGND VGND VPWR VPWR dadda_fa_1_69_6/B
+ dadda_fa_1_68_8/A sky130_fd_sc_hd__fa_1
XTAP_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_45_1 dadda_fa_3_45_1/A dadda_fa_3_45_1/B dadda_fa_3_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_0/CIN dadda_fa_4_45_2/A sky130_fd_sc_hd__fa_1
XTAP_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_22_0 dadda_fa_6_22_0/A dadda_fa_6_22_0/B dadda_fa_6_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_23_0/B dadda_fa_7_22_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_38_0 dadda_fa_3_38_0/A dadda_fa_3_38_0/B dadda_fa_3_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_0/B dadda_fa_4_38_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$730 U$$730/A U$$796/B VGND VGND VPWR VPWR U$$730/X sky130_fd_sc_hd__xor2_1
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_666_ _674_/CLK _666_/D VGND VGND VPWR VPWR _666_/Q sky130_fd_sc_hd__dfxtp_1
XU$$741 U$$878/A1 U$$747/A2 U$$880/A1 U$$747/B2 VGND VGND VPWR VPWR U$$742/A sky130_fd_sc_hd__a22o_1
XFILLER_189_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$752 U$$752/A U$$804/B VGND VGND VPWR VPWR U$$752/X sky130_fd_sc_hd__xor2_1
XFILLER_1_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$763 U$$900/A1 U$$765/A2 U$$900/B1 U$$765/B2 VGND VGND VPWR VPWR U$$764/A sky130_fd_sc_hd__a22o_1
XFILLER_204_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$774 U$$774/A U$$816/B VGND VGND VPWR VPWR U$$774/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_597_ _598_/CLK _597_/D VGND VGND VPWR VPWR _597_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$785 U$$922/A1 U$$819/A2 U$$785/B1 U$$819/B2 VGND VGND VPWR VPWR U$$786/A sky130_fd_sc_hd__a22o_1
XU$$796 U$$796/A U$$796/B VGND VGND VPWR VPWR U$$796/X sky130_fd_sc_hd__xor2_1
XFILLER_90_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_2 _456_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_97_4 U$$3925/X U$$4058/X U$$4191/X VGND VGND VPWR VPWR dadda_fa_3_98_1/CIN
+ dadda_fa_3_97_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1630 U$$985/A1 VGND VGND VPWR VPWR U$$435/B1 sky130_fd_sc_hd__buf_6
XFILLER_67_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1641 U$$3584/B1 VGND VGND VPWR VPWR U$$24/A1 sky130_fd_sc_hd__buf_4
XFILLER_99_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1652 U$$4404/B1 VGND VGND VPWR VPWR U$$4269/A1 sky130_fd_sc_hd__buf_6
XFILLER_141_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1663 U$$2895/A1 VGND VGND VPWR VPWR U$$18/A1 sky130_fd_sc_hd__buf_6
XFILLER_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1674 U$$2756/A1 VGND VGND VPWR VPWR U$$838/A1 sky130_fd_sc_hd__buf_4
XFILLER_153_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1685 U$$4259/B1 VGND VGND VPWR VPWR U$$3713/A1 sky130_fd_sc_hd__buf_8
XFILLER_154_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1696 U$$556/B1 VGND VGND VPWR VPWR U$$695/A1 sky130_fd_sc_hd__buf_6
XFILLER_141_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_478 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_40_0 U$$1550/X U$$1683/X U$$1816/X VGND VGND VPWR VPWR dadda_fa_3_41_0/B
+ dadda_fa_3_40_2/B sky130_fd_sc_hd__fa_1
XFILLER_26_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2170 U$$2170/A U$$2170/B VGND VGND VPWR VPWR U$$2170/X sky130_fd_sc_hd__xor2_1
XU$$2181 U$$2866/A1 U$$2185/A2 U$$2318/B1 U$$2185/B2 VGND VGND VPWR VPWR U$$2182/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2192 _647_/Q VGND VGND VPWR VPWR U$$2192/Y sky130_fd_sc_hd__inv_1
XFILLER_50_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1480 U$$658/A1 U$$1486/A2 U$$384/B1 U$$1486/B2 VGND VGND VPWR VPWR U$$1481/A sky130_fd_sc_hd__a22o_1
XU$$1491 U$$1491/A U$$1501/B VGND VGND VPWR VPWR U$$1491/X sky130_fd_sc_hd__xor2_1
XFILLER_210_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1092 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_2 U$$2305/X U$$2438/X U$$2571/X VGND VGND VPWR VPWR dadda_fa_2_86_3/A
+ dadda_fa_2_85_5/A sky130_fd_sc_hd__fa_1
XFILLER_131_431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_62_1 dadda_fa_4_62_1/A dadda_fa_4_62_1/B dadda_fa_4_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/B dadda_fa_5_62_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_78_1 U$$1626/X U$$1759/X U$$1892/X VGND VGND VPWR VPWR dadda_fa_2_79_0/CIN
+ dadda_fa_2_78_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_55_0 dadda_fa_4_55_0/A dadda_fa_4_55_0/B dadda_fa_4_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/A dadda_fa_5_55_1/A sky130_fd_sc_hd__fa_1
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$110 _534_/Q _406_/Q VGND VGND VPWR VPWR final_adder.U$$605/B1 final_adder.U$$732/A
+ sky130_fd_sc_hd__ha_2
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$121 _545_/Q _417_/Q VGND VGND VPWR VPWR final_adder.U$$249/B1 final_adder.U$$743/A
+ sky130_fd_sc_hd__ha_2
XFILLER_100_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$132 final_adder.U$$627/A final_adder.U$$626/A VGND VGND VPWR VPWR
+ final_adder.U$$258/B sky130_fd_sc_hd__and2_1
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$143 final_adder.U$$637/A final_adder.U$$509/B1 final_adder.U$$143/B1
+ VGND VGND VPWR VPWR final_adder.U$$143/X sky130_fd_sc_hd__a21o_1
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$154 final_adder.U$$649/A final_adder.U$$648/A VGND VGND VPWR VPWR
+ final_adder.U$$268/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$165 final_adder.U$$659/A final_adder.U$$531/B1 final_adder.U$$165/B1
+ VGND VGND VPWR VPWR final_adder.U$$165/X sky130_fd_sc_hd__a21o_1
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$176 final_adder.U$$671/A final_adder.U$$670/A VGND VGND VPWR VPWR
+ final_adder.U$$280/B sky130_fd_sc_hd__and2_1
X_520_ _520_/CLK _520_/D VGND VGND VPWR VPWR _520_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$187 final_adder.U$$681/A final_adder.U$$553/B1 final_adder.U$$187/B1
+ VGND VGND VPWR VPWR final_adder.U$$187/X sky130_fd_sc_hd__a21o_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater391 U$$963/X VGND VGND VPWR VPWR U$$1093/A2 sky130_fd_sc_hd__buf_6
XFILLER_57_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$198 final_adder.U$$693/A final_adder.U$$692/A VGND VGND VPWR VPWR
+ final_adder.U$$290/A sky130_fd_sc_hd__and2_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_451_ _451_/CLK _451_/D VGND VGND VPWR VPWR _451_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_382_ _560_/CLK _382_/D VGND VGND VPWR VPWR _382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_74_2 U$$1485/X U$$1618/X VGND VGND VPWR VPWR dadda_fa_1_75_8/B dadda_fa_2_74_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_107_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_73_0 U$$684/Y U$$818/X U$$951/X VGND VGND VPWR VPWR dadda_fa_1_74_7/B
+ dadda_fa_1_73_8/B sky130_fd_sc_hd__fa_1
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput150 c[119] VGND VGND VPWR VPWR input150/X sky130_fd_sc_hd__dlymetal6s2s_1
XU$$134_1716 VGND VGND VPWR VPWR U$$134_1716/HI U$$134/B1 sky130_fd_sc_hd__conb_1
XFILLER_76_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput161 c[13] VGND VGND VPWR VPWR input161/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_551 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput172 c[23] VGND VGND VPWR VPWR input172/X sky130_fd_sc_hd__buf_2
XFILLER_3_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput183 c[33] VGND VGND VPWR VPWR input183/X sky130_fd_sc_hd__clkbuf_4
Xinput194 c[43] VGND VGND VPWR VPWR input194/X sky130_fd_sc_hd__clkbuf_1
XTAP_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_649_ _660_/CLK _649_/D VGND VGND VPWR VPWR _649_/Q sky130_fd_sc_hd__dfxtp_2
XU$$560 U$$695/B1 U$$574/A2 U$$562/A1 U$$574/B2 VGND VGND VPWR VPWR U$$561/A sky130_fd_sc_hd__a22o_1
XFILLER_17_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$571 U$$571/A U$$589/B VGND VGND VPWR VPWR U$$571/X sky130_fd_sc_hd__xor2_1
XU$$582 U$$582/A1 U$$616/A2 U$$582/B1 U$$616/B2 VGND VGND VPWR VPWR U$$583/A sky130_fd_sc_hd__a22o_1
XFILLER_204_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$593 U$$593/A U$$665/B VGND VGND VPWR VPWR U$$593/X sky130_fd_sc_hd__xor2_1
XFILLER_32_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_95_1 U$$2990/X U$$3123/X U$$3256/X VGND VGND VPWR VPWR dadda_fa_3_96_0/CIN
+ dadda_fa_3_95_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_145_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_72_0 dadda_fa_5_72_0/A dadda_fa_5_72_0/B dadda_fa_5_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_73_0/A dadda_fa_6_72_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1460 U$$4450/B1 VGND VGND VPWR VPWR U$$68/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_88_0 U$$3508/X U$$3641/X U$$3774/X VGND VGND VPWR VPWR dadda_fa_3_89_0/B
+ dadda_fa_3_88_2/B sky130_fd_sc_hd__fa_1
XFILLER_132_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1471 U$$3902/A1 VGND VGND VPWR VPWR U$$66/A1 sky130_fd_sc_hd__buf_4
Xrepeater1482 _580_/Q VGND VGND VPWR VPWR U$$4446/B1 sky130_fd_sc_hd__buf_6
XFILLER_98_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1493 U$$3485/A1 VGND VGND VPWR VPWR U$$745/A1 sky130_fd_sc_hd__buf_4
XU$$3285_1748 VGND VGND VPWR VPWR U$$3285_1748/HI U$$3285/B1 sky130_fd_sc_hd__conb_1
XFILLER_67_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_71_8 dadda_fa_1_71_8/A dadda_fa_1_71_8/B dadda_fa_1_71_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_72_3/A dadda_fa_3_71_0/A sky130_fd_sc_hd__fa_2
XFILLER_141_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_64_7 dadda_fa_1_64_7/A dadda_fa_1_64_7/B dadda_fa_1_64_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_2/CIN dadda_fa_2_64_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_57_6 U$$3579/X U$$3712/X U$$3845/X VGND VGND VPWR VPWR dadda_fa_2_58_2/B
+ dadda_fa_2_57_5/B sky130_fd_sc_hd__fa_1
XFILLER_41_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4387_1770 VGND VGND VPWR VPWR U$$4387_1770/HI U$$4387/A sky130_fd_sc_hd__conb_1
XFILLER_55_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_9_0 dadda_fa_7_9_0/A dadda_fa_7_9_0/B dadda_fa_7_9_0/CIN VGND VGND VPWR
+ VPWR _434_/D _305_/D sky130_fd_sc_hd__fa_1
XU$$4461_1809 VGND VGND VPWR VPWR U$$4461_1809/HI U$$4461/B sky130_fd_sc_hd__conb_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_87_0 dadda_fa_7_87_0/A dadda_fa_7_87_0/B dadda_fa_7_87_0/CIN VGND VGND
+ VPWR VPWR _512_/D _383_/D sky130_fd_sc_hd__fa_1
XFILLER_202_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_90_0 dadda_fa_1_90_0/A U$$1916/X U$$2049/X VGND VGND VPWR VPWR dadda_fa_2_91_4/A
+ dadda_fa_2_90_5/A sky130_fd_sc_hd__fa_1
XFILLER_105_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4308 U$$4308/A _679_/Q VGND VGND VPWR VPWR U$$4308/X sky130_fd_sc_hd__xor2_1
XU$$4319 _584_/Q U$$4327/A2 _585_/Q U$$4319/B2 VGND VGND VPWR VPWR U$$4320/A sky130_fd_sc_hd__a22o_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3607 U$$3607/A U$$3609/B VGND VGND VPWR VPWR U$$3607/X sky130_fd_sc_hd__xor2_1
XU$$3618 U$$3618/A1 U$$3662/A2 _577_/Q U$$3662/B2 VGND VGND VPWR VPWR U$$3619/A sky130_fd_sc_hd__a22o_1
XFILLER_92_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3629 U$$3629/A U$$3675/B VGND VGND VPWR VPWR U$$3629/X sky130_fd_sc_hd__xor2_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_102_0 dadda_fa_6_102_0/A dadda_fa_6_102_0/B dadda_fa_6_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_103_0/B dadda_fa_7_102_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2906 U$$2906/A U$$2988/B VGND VGND VPWR VPWR U$$2906/X sky130_fd_sc_hd__xor2_1
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 _185_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2917 U$$999/A1 U$$2943/A2 U$$3193/A1 U$$2943/B2 VGND VGND VPWR VPWR U$$2918/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2928 U$$2928/A U$$2928/B VGND VGND VPWR VPWR U$$2928/X sky130_fd_sc_hd__xor2_1
XANTENNA_211 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_503_ _503_/CLK _503_/D VGND VGND VPWR VPWR _503_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2939 U$$4035/A1 U$$2973/A2 U$$4035/B1 U$$2973/B2 VGND VGND VPWR VPWR U$$2940/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_22_3 U$$1514/X U$$1558/B input171/X VGND VGND VPWR VPWR dadda_fa_4_23_1/B
+ dadda_fa_4_22_2/CIN sky130_fd_sc_hd__fa_1
XANTENNA_233 _188_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 _193_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_255 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_266 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_434_ _435_/CLK _434_/D VGND VGND VPWR VPWR _434_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_277 _212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_288 _214_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_299 _234_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_365_ _494_/CLK _365_/D VGND VGND VPWR VPWR _365_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_296_ _431_/CLK _296_/D VGND VGND VPWR VPWR _296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_clk _616_/CLK VGND VGND VPWR VPWR _488_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_67_5 dadda_fa_2_67_5/A dadda_fa_2_67_5/B dadda_fa_2_67_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_2/A dadda_fa_4_67_0/A sky130_fd_sc_hd__fa_1
XFILLER_122_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$390 U$$527/A1 U$$392/A2 U$$392/A1 U$$392/B2 VGND VGND VPWR VPWR U$$391/A sky130_fd_sc_hd__a22o_1
XFILLER_33_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4419_1788 VGND VGND VPWR VPWR U$$4419_1788/HI U$$4419/B sky130_fd_sc_hd__conb_1
XFILLER_160_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1290 U$$382/B1 VGND VGND VPWR VPWR U$$658/A1 sky130_fd_sc_hd__buf_6
XFILLER_99_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_62_4 U$$3988/X U$$4121/X U$$4254/X VGND VGND VPWR VPWR dadda_fa_2_63_1/CIN
+ dadda_fa_2_62_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_55_3 U$$1979/X U$$2112/X U$$2245/X VGND VGND VPWR VPWR dadda_fa_2_56_1/B
+ dadda_fa_2_55_4/B sky130_fd_sc_hd__fa_1
XFILLER_80_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_32_2 dadda_fa_4_32_2/A dadda_fa_4_32_2/B dadda_fa_4_32_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/CIN dadda_fa_5_32_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_48_2 U$$901/X U$$1034/X U$$1167/X VGND VGND VPWR VPWR dadda_fa_2_49_1/CIN
+ dadda_fa_2_48_4/B sky130_fd_sc_hd__fa_1
XFILLER_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_25_1 dadda_fa_4_25_1/A dadda_fa_4_25_1/B dadda_fa_4_25_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/B dadda_fa_5_25_1/B sky130_fd_sc_hd__fa_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_18_0 U$$1107/X U$$1240/X U$$1288/B VGND VGND VPWR VPWR dadda_fa_5_19_0/A
+ dadda_fa_5_18_1/A sky130_fd_sc_hd__fa_1
XFILLER_208_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_751 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4105 U$$4105/A1 U$$4107/A2 U$$4105/B1 U$$4105/B2 VGND VGND VPWR VPWR U$$4106/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4116 U$$4116/A1 U$$4140/A2 U$$4392/A1 U$$4140/B2 VGND VGND VPWR VPWR U$$4117/A
+ sky130_fd_sc_hd__a22o_1
XU$$4127 U$$4127/A U$$4141/B VGND VGND VPWR VPWR U$$4127/X sky130_fd_sc_hd__xor2_1
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4138 U$$4273/B1 U$$4140/A2 U$$4140/A1 U$$4140/B2 VGND VGND VPWR VPWR U$$4139/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4149 U$$4149/A U$$4183/B VGND VGND VPWR VPWR U$$4149/X sky130_fd_sc_hd__xor2_1
XFILLER_101_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3404 U$$3404/A1 U$$3404/A2 U$$4502/A1 U$$3404/B2 VGND VGND VPWR VPWR U$$3405/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3415 U$$3415/A U$$3423/B VGND VGND VPWR VPWR U$$3415/X sky130_fd_sc_hd__xor2_1
XU$$3426 _666_/Q VGND VGND VPWR VPWR U$$3428/B sky130_fd_sc_hd__inv_1
XU$$3437 U$$3437/A1 U$$3479/A2 U$$3713/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3438/A
+ sky130_fd_sc_hd__a22o_1
XU$$4483_1820 VGND VGND VPWR VPWR U$$4483_1820/HI U$$4483/B sky130_fd_sc_hd__conb_1
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2703 U$$2838/B1 U$$2705/A2 U$$2705/A1 U$$2705/B2 VGND VGND VPWR VPWR U$$2704/A
+ sky130_fd_sc_hd__a22o_1
XU$$3448 U$$3448/A U$$3498/B VGND VGND VPWR VPWR U$$3448/X sky130_fd_sc_hd__xor2_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2714 U$$2714/A U$$2734/B VGND VGND VPWR VPWR U$$2714/X sky130_fd_sc_hd__xor2_1
XFILLER_46_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3459 U$$4007/A1 U$$3559/A2 U$$3735/A1 U$$3559/B2 VGND VGND VPWR VPWR U$$3460/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2725 U$$2725/A1 U$$2729/A2 _610_/Q U$$2729/B2 VGND VGND VPWR VPWR U$$2726/A sky130_fd_sc_hd__a22o_1
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2736 U$$2736/A U$$2739/A VGND VGND VPWR VPWR U$$2736/X sky130_fd_sc_hd__xor2_1
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2747 U$$2747/A U$$2787/B VGND VGND VPWR VPWR U$$2747/X sky130_fd_sc_hd__xor2_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2758 U$$2893/B1 U$$2788/A2 U$$3717/B1 U$$2788/B2 VGND VGND VPWR VPWR U$$2759/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_0 U$$47/X U$$180/X U$$313/X VGND VGND VPWR VPWR dadda_fa_4_21_0/B dadda_fa_4_20_1/CIN
+ sky130_fd_sc_hd__fa_1
XU$$2769 U$$2769/A U$$2827/B VGND VGND VPWR VPWR U$$2769/X sky130_fd_sc_hd__xor2_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_417_ _547_/CLK _417_/D VGND VGND VPWR VPWR _417_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_348_ _476_/CLK _348_/D VGND VGND VPWR VPWR _348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_279_ _523_/CLK _279_/D VGND VGND VPWR VPWR _279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_72_3 dadda_fa_2_72_3/A dadda_fa_2_72_3/B dadda_fa_2_72_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/B dadda_fa_3_72_3/B sky130_fd_sc_hd__fa_1
XFILLER_29_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_65_2 dadda_fa_2_65_2/A dadda_fa_2_65_2/B dadda_fa_2_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/A dadda_fa_3_65_3/A sky130_fd_sc_hd__fa_1
XFILLER_9_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater902 U$$4389/X VGND VGND VPWR VPWR U$$4496/B2 sky130_fd_sc_hd__buf_4
XFILLER_69_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$709 final_adder.U$$709/A final_adder.U$$709/B VGND VGND VPWR VPWR
+ _255_/D sky130_fd_sc_hd__xor2_1
Xrepeater913 U$$4203/B VGND VGND VPWR VPWR U$$4197/B sky130_fd_sc_hd__buf_6
XFILLER_64_1099 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_42_1 dadda_fa_5_42_1/A dadda_fa_5_42_1/B dadda_fa_5_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_43_0/B dadda_fa_7_42_0/A sky130_fd_sc_hd__fa_2
Xrepeater924 U$$4084/B VGND VGND VPWR VPWR U$$4096/B sky130_fd_sc_hd__buf_6
Xrepeater935 U$$3943/B VGND VGND VPWR VPWR U$$3949/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_58_1 dadda_fa_2_58_1/A dadda_fa_2_58_1/B dadda_fa_2_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_0/CIN dadda_fa_3_58_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater946 U$$3836/A VGND VGND VPWR VPWR U$$3835/A sky130_fd_sc_hd__buf_6
Xrepeater957 U$$3556/B VGND VGND VPWR VPWR U$$3561/A sky130_fd_sc_hd__buf_6
Xdadda_fa_5_35_0 dadda_fa_5_35_0/A dadda_fa_5_35_0/B dadda_fa_5_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_36_0/A dadda_fa_6_35_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater968 U$$3363/B VGND VGND VPWR VPWR U$$3343/B sky130_fd_sc_hd__buf_12
XFILLER_110_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater979 U$$3286/B VGND VGND VPWR VPWR U$$3208/B sky130_fd_sc_hd__buf_6
XFILLER_209_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3960 U$$4369/B1 U$$3970/A2 U$$4236/A1 U$$3970/B2 VGND VGND VPWR VPWR U$$3961/A
+ sky130_fd_sc_hd__a22o_1
XU$$3971 U$$3971/A U$$3973/A VGND VGND VPWR VPWR U$$3971/X sky130_fd_sc_hd__xor2_1
XFILLER_24_215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3982 U$$3982/A U$$4036/B VGND VGND VPWR VPWR U$$3982/X sky130_fd_sc_hd__xor2_1
XU$$3993 U$$4402/B1 U$$4005/A2 U$$4269/A1 U$$4005/B2 VGND VGND VPWR VPWR U$$3994/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1915_1726 VGND VGND VPWR VPWR U$$1915_1726/HI U$$1915/B1 sky130_fd_sc_hd__conb_1
XFILLER_75_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput262 _272_/Q VGND VGND VPWR VPWR o[104] sky130_fd_sc_hd__buf_2
XFILLER_160_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput273 _282_/Q VGND VGND VPWR VPWR o[114] sky130_fd_sc_hd__buf_2
XFILLER_161_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput284 _292_/Q VGND VGND VPWR VPWR o[124] sky130_fd_sc_hd__buf_2
XFILLER_82_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput295 _187_/Q VGND VGND VPWR VPWR o[19] sky130_fd_sc_hd__buf_2
XFILLER_102_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_60_1 U$$2388/X U$$2521/X U$$2654/X VGND VGND VPWR VPWR dadda_fa_2_61_0/CIN
+ dadda_fa_2_60_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_53_0 U$$379/X U$$512/X U$$645/X VGND VGND VPWR VPWR dadda_fa_2_54_0/B
+ dadda_fa_2_53_3/B sky130_fd_sc_hd__fa_1
XFILLER_68_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1309 U$$76/A1 U$$1309/A2 U$$78/A1 U$$1309/B2 VGND VGND VPWR VPWR U$$1310/A sky130_fd_sc_hd__a22o_1
XFILLER_43_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_202_ _213_/CLK _202_/D VGND VGND VPWR VPWR _202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_927 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$280_1741 VGND VGND VPWR VPWR U$$280_1741/HI U$$280/A1 sky130_fd_sc_hd__conb_1
XFILLER_211_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4107_1762 VGND VGND VPWR VPWR U$$4107_1762/HI U$$4107/B1 sky130_fd_sc_hd__conb_1
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_82_2 dadda_fa_3_82_2/A dadda_fa_3_82_2/B dadda_fa_3_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_1/A dadda_fa_4_82_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_3_75_1 dadda_fa_3_75_1/A dadda_fa_3_75_1/B dadda_fa_3_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_0/CIN dadda_fa_4_75_2/A sky130_fd_sc_hd__fa_1
XFILLER_151_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_52_0 dadda_fa_6_52_0/A dadda_fa_6_52_0/B dadda_fa_6_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_53_0/B dadda_fa_7_52_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_68_0 dadda_fa_3_68_0/A dadda_fa_3_68_0/B dadda_fa_3_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_0/B dadda_fa_4_68_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3201 U$$4434/A1 U$$3235/A2 U$$4436/A1 U$$3235/B2 VGND VGND VPWR VPWR U$$3202/A
+ sky130_fd_sc_hd__a22o_1
XU$$3212 U$$3212/A U$$3232/B VGND VGND VPWR VPWR U$$3212/X sky130_fd_sc_hd__xor2_1
XFILLER_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3223 U$$4317/B1 U$$3231/A2 U$$4184/A1 U$$3231/B2 VGND VGND VPWR VPWR U$$3224/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_150_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_111_2 dadda_fa_4_111_2/A dadda_fa_4_111_2/B dadda_fa_4_111_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_112_0/CIN dadda_fa_5_111_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$16 _440_/Q _312_/Q VGND VGND VPWR VPWR final_adder.U$$511/B1 final_adder.U$$638/A
+ sky130_fd_sc_hd__ha_2
XFILLER_47_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3234 U$$3234/A U$$3276/B VGND VGND VPWR VPWR U$$3234/X sky130_fd_sc_hd__xor2_1
XFILLER_93_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2500 U$$2909/B1 U$$2550/A2 U$$2774/B1 U$$2550/B2 VGND VGND VPWR VPWR U$$2501/A
+ sky130_fd_sc_hd__a22o_1
XU$$3245 U$$4065/B1 U$$3283/A2 U$$3245/B1 U$$3283/B2 VGND VGND VPWR VPWR U$$3246/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3256 U$$3256/A U$$3256/B VGND VGND VPWR VPWR U$$3256/X sky130_fd_sc_hd__xor2_1
XU$$2511 U$$2511/A U$$2551/B VGND VGND VPWR VPWR U$$2511/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$27 _451_/Q _323_/Q VGND VGND VPWR VPWR final_adder.U$$155/B1 final_adder.U$$649/A
+ sky130_fd_sc_hd__ha_2
XFILLER_94_1004 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$38 _462_/Q _334_/Q VGND VGND VPWR VPWR final_adder.U$$533/B1 final_adder.U$$660/A
+ sky130_fd_sc_hd__ha_1
XU$$3267 _606_/Q U$$3273/A2 U$$3952/B1 U$$3273/B2 VGND VGND VPWR VPWR U$$3268/A sky130_fd_sc_hd__a22o_1
XFILLER_4_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2522 U$$56/A1 U$$2524/A2 U$$2796/B1 U$$2524/B2 VGND VGND VPWR VPWR U$$2523/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_104_1 dadda_fa_4_104_1/A dadda_fa_4_104_1/B dadda_fa_4_104_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/B dadda_fa_5_104_1/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$49 _473_/Q _345_/Q VGND VGND VPWR VPWR final_adder.U$$177/B1 final_adder.U$$671/A
+ sky130_fd_sc_hd__ha_1
XU$$2533 U$$2533/A _653_/Q VGND VGND VPWR VPWR U$$2533/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3278 U$$3278/A U$$3288/A VGND VGND VPWR VPWR U$$3278/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3289 _664_/Q VGND VGND VPWR VPWR U$$3291/B sky130_fd_sc_hd__inv_1
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2544 U$$3229/A1 U$$2566/A2 U$$628/A1 U$$2566/B2 VGND VGND VPWR VPWR U$$2545/A
+ sky130_fd_sc_hd__a22o_1
XU$$2555 U$$2555/A U$$2597/B VGND VGND VPWR VPWR U$$2555/X sky130_fd_sc_hd__xor2_1
XU$$1810 U$$1810/A U$$1852/B VGND VGND VPWR VPWR U$$1810/X sky130_fd_sc_hd__xor2_1
XFILLER_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1821 U$$3054/A1 U$$1785/X U$$3193/A1 U$$1786/X VGND VGND VPWR VPWR U$$1822/A sky130_fd_sc_hd__a22o_1
XU$$2566 U$$922/A1 U$$2566/A2 U$$924/A1 U$$2566/B2 VGND VGND VPWR VPWR U$$2567/A sky130_fd_sc_hd__a22o_1
XFILLER_179_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1832 U$$1832/A U$$1852/B VGND VGND VPWR VPWR U$$1832/X sky130_fd_sc_hd__xor2_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2577 U$$2577/A U$$2583/B VGND VGND VPWR VPWR U$$2577/X sky130_fd_sc_hd__xor2_1
XU$$1843 U$$1843/A1 U$$1843/A2 U$$3352/A1 U$$1843/B2 VGND VGND VPWR VPWR U$$1844/A
+ sky130_fd_sc_hd__a22o_1
XU$$2588 U$$2725/A1 U$$2588/A2 U$$2588/B1 U$$2588/B2 VGND VGND VPWR VPWR U$$2589/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1854 U$$1854/A U$$1884/B VGND VGND VPWR VPWR U$$1854/X sky130_fd_sc_hd__xor2_1
XU$$2599 U$$2599/A U$$2603/A VGND VGND VPWR VPWR U$$2599/X sky130_fd_sc_hd__xor2_1
XFILLER_15_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1865 U$$358/A1 U$$1785/X U$$86/A1 U$$1786/X VGND VGND VPWR VPWR U$$1866/A sky130_fd_sc_hd__a22o_1
XU$$1876 U$$1876/A U$$1916/B VGND VGND VPWR VPWR U$$1876/X sky130_fd_sc_hd__xor2_1
XU$$1887 U$$3255/B1 U$$1897/A2 U$$3122/A1 U$$1897/B2 VGND VGND VPWR VPWR U$$1888/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1898 U$$1898/A U$$1917/A VGND VGND VPWR VPWR U$$1898/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_125_0 dadda_fa_7_125_0/A dadda_fa_7_125_0/B dadda_fa_7_125_0/CIN VGND
+ VGND VPWR VPWR _550_/D _421_/D sky130_fd_sc_hd__fa_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_774 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1043 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_992 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_985 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_70_0 dadda_fa_2_70_0/A dadda_fa_2_70_0/B dadda_fa_2_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_0/B dadda_fa_3_70_2/B sky130_fd_sc_hd__fa_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater710 U$$3769/B2 VGND VGND VPWR VPWR U$$3743/B2 sky130_fd_sc_hd__buf_6
XFILLER_97_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater721 U$$3688/B2 VGND VGND VPWR VPWR U$$3696/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$517 final_adder.U$$644/A final_adder.U$$644/B final_adder.U$$517/B1
+ VGND VGND VPWR VPWR final_adder.U$$645/B sky130_fd_sc_hd__a21o_1
XFILLER_111_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater732 U$$3555/B2 VGND VGND VPWR VPWR U$$3545/B2 sky130_fd_sc_hd__buf_4
XFILLER_57_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$539 final_adder.U$$666/A final_adder.U$$666/B final_adder.U$$539/B1
+ VGND VGND VPWR VPWR final_adder.U$$667/B sky130_fd_sc_hd__a21o_1
XFILLER_96_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater743 U$$3285/B2 VGND VGND VPWR VPWR U$$3235/B2 sky130_fd_sc_hd__buf_6
Xrepeater754 U$$3148/B2 VGND VGND VPWR VPWR U$$3110/B2 sky130_fd_sc_hd__buf_8
Xrepeater765 U$$2882/X VGND VGND VPWR VPWR U$$3005/B2 sky130_fd_sc_hd__buf_4
Xrepeater776 U$$2832/B2 VGND VGND VPWR VPWR U$$2812/B2 sky130_fd_sc_hd__buf_6
Xrepeater787 U$$2729/B2 VGND VGND VPWR VPWR U$$2687/B2 sky130_fd_sc_hd__buf_4
XU$$4480 U$$4480/A1 U$$4388/X U$$4482/A1 U$$4480/B2 VGND VGND VPWR VPWR U$$4481/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater798 U$$2471/X VGND VGND VPWR VPWR U$$2580/B2 sky130_fd_sc_hd__buf_6
XU$$4491 U$$4491/A U$$4491/B VGND VGND VPWR VPWR U$$4491/X sky130_fd_sc_hd__xor2_1
XFILLER_37_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_91_clk _628_/CLK VGND VGND VPWR VPWR _541_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$3790 U$$3790/A U$$3804/B VGND VGND VPWR VPWR U$$3790/X sky130_fd_sc_hd__xor2_1
XFILLER_198_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_724 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_92_1 dadda_fa_4_92_1/A dadda_fa_4_92_1/B dadda_fa_4_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/B dadda_fa_5_92_1/B sky130_fd_sc_hd__fa_1
Xclkbuf_3_0__f_clk clkbuf_2_0_0_clk/X VGND VGND VPWR VPWR _442_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_85_0 dadda_fa_4_85_0/A dadda_fa_4_85_0/B dadda_fa_4_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/A dadda_fa_5_85_1/A sky130_fd_sc_hd__fa_1
XFILLER_107_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_106_3 dadda_fa_3_106_3/A dadda_fa_3_106_3/B dadda_fa_3_106_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_107_1/B dadda_fa_4_106_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3011_1744 VGND VGND VPWR VPWR U$$3011_1744/HI U$$3011/B1 sky130_fd_sc_hd__conb_1
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$901 U$$901/A U$$907/B VGND VGND VPWR VPWR U$$901/X sky130_fd_sc_hd__xor2_1
XU$$912 U$$912/A1 U$$956/A2 U$$912/B1 U$$956/B2 VGND VGND VPWR VPWR U$$913/A sky130_fd_sc_hd__a22o_1
XFILLER_28_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$923 U$$923/A U$$925/B VGND VGND VPWR VPWR U$$923/X sky130_fd_sc_hd__xor2_1
XFILLER_90_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$934 U$$934/A1 U$$826/X U$$936/A1 U$$827/X VGND VGND VPWR VPWR U$$935/A sky130_fd_sc_hd__a22o_1
XFILLER_204_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$945 U$$945/A U$$951/B VGND VGND VPWR VPWR U$$945/X sky130_fd_sc_hd__xor2_1
XU$$956 U$$956/A1 U$$956/A2 U$$956/B1 U$$956/B2 VGND VGND VPWR VPWR U$$957/A sky130_fd_sc_hd__a22o_1
XFILLER_189_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$967 U$$967/A1 U$$995/A2 U$$969/A1 U$$995/B2 VGND VGND VPWR VPWR U$$968/A sky130_fd_sc_hd__a22o_1
XU$$1106 U$$969/A1 U$$1150/A2 U$$971/A1 U$$1150/B2 VGND VGND VPWR VPWR U$$1107/A sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_82_clk _628_/CLK VGND VGND VPWR VPWR _660_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$978 U$$978/A U$$980/B VGND VGND VPWR VPWR U$$978/X sky130_fd_sc_hd__xor2_1
XU$$1117 U$$1117/A U$$1151/B VGND VGND VPWR VPWR U$$1117/X sky130_fd_sc_hd__xor2_1
XFILLER_203_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1128 U$$991/A1 U$$1194/A2 U$$993/A1 U$$1194/B2 VGND VGND VPWR VPWR U$$1129/A sky130_fd_sc_hd__a22o_1
XU$$989 U$$989/A1 U$$995/A2 U$$32/A1 U$$995/B2 VGND VGND VPWR VPWR U$$990/A sky130_fd_sc_hd__a22o_1
XFILLER_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1139 U$$1139/A U$$1147/B VGND VGND VPWR VPWR U$$1139/X sky130_fd_sc_hd__xor2_1
XFILLER_31_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1010 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1040 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_831 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_42_4 dadda_fa_2_42_4/A dadda_fa_2_42_4/B dadda_fa_2_42_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_43_1/CIN dadda_fa_3_42_3/CIN sky130_fd_sc_hd__fa_1
XU$$3020 U$$3020/A1 U$$3054/A2 U$$3157/B1 U$$3054/B2 VGND VGND VPWR VPWR U$$3021/A
+ sky130_fd_sc_hd__a22o_1
XU$$3031 U$$3031/A U$$3049/B VGND VGND VPWR VPWR U$$3031/X sky130_fd_sc_hd__xor2_1
XFILLER_53_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3042 U$$3042/A1 U$$3082/A2 U$$3042/B1 U$$3082/B2 VGND VGND VPWR VPWR U$$3043/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_35_3 U$$1540/X U$$1673/X U$$1806/X VGND VGND VPWR VPWR dadda_fa_3_36_1/B
+ dadda_fa_3_35_3/B sky130_fd_sc_hd__fa_1
XU$$3053 U$$3053/A U$$3077/B VGND VGND VPWR VPWR U$$3053/X sky130_fd_sc_hd__xor2_1
XFILLER_81_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3064 U$$4434/A1 U$$3066/A2 U$$4436/A1 U$$3066/B2 VGND VGND VPWR VPWR U$$3065/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2330 _650_/Q VGND VGND VPWR VPWR U$$2332/B sky130_fd_sc_hd__inv_1
XU$$3075 U$$3075/A U$$3077/B VGND VGND VPWR VPWR U$$3075/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_73_clk _634_/CLK VGND VGND VPWR VPWR _514_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$3086 U$$3221/B1 U$$3120/A2 U$$3088/A1 U$$3120/B2 VGND VGND VPWR VPWR U$$3087/A
+ sky130_fd_sc_hd__a22o_1
XU$$2341 U$$2478/A1 U$$2367/A2 U$$2343/A1 U$$2367/B2 VGND VGND VPWR VPWR U$$2342/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2352 U$$2352/A U$$2400/B VGND VGND VPWR VPWR U$$2352/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_28_2 U$$861/X U$$994/X U$$1127/X VGND VGND VPWR VPWR dadda_fa_3_29_2/B
+ dadda_fa_3_28_3/CIN sky130_fd_sc_hd__fa_1
XU$$3097 U$$3097/A U$$3111/B VGND VGND VPWR VPWR U$$3097/X sky130_fd_sc_hd__xor2_1
XU$$2363 U$$3046/B1 U$$2387/A2 U$$582/B1 U$$2387/B2 VGND VGND VPWR VPWR U$$2364/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2374 U$$2374/A U$$2418/B VGND VGND VPWR VPWR U$$2374/X sky130_fd_sc_hd__xor2_1
XFILLER_179_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1640 U$$1640/A _639_/Q VGND VGND VPWR VPWR U$$1640/X sky130_fd_sc_hd__xor2_1
XU$$2385 U$$4027/B1 U$$2387/A2 U$$467/B1 U$$2387/B2 VGND VGND VPWR VPWR U$$2386/A
+ sky130_fd_sc_hd__a22o_1
XU$$2396 U$$2396/A U$$2400/B VGND VGND VPWR VPWR U$$2396/X sky130_fd_sc_hd__xor2_1
XU$$1651 U$$1651/A U$$1723/B VGND VGND VPWR VPWR U$$1651/X sky130_fd_sc_hd__xor2_1
XU$$1662 U$$840/A1 U$$1684/A2 U$$840/B1 U$$1684/B2 VGND VGND VPWR VPWR U$$1663/A sky130_fd_sc_hd__a22o_1
XU$$1673 U$$1673/A U$$1711/B VGND VGND VPWR VPWR U$$1673/X sky130_fd_sc_hd__xor2_1
XFILLER_201_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1684 U$$3054/A1 U$$1684/A2 U$$42/A1 U$$1684/B2 VGND VGND VPWR VPWR U$$1685/A sky130_fd_sc_hd__a22o_1
XFILLER_72_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1695 U$$1695/A U$$1723/B VGND VGND VPWR VPWR U$$1695/X sky130_fd_sc_hd__xor2_1
XFILLER_72_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$303 final_adder.U$$302/A final_adder.U$$221/X final_adder.U$$223/X
+ VGND VGND VPWR VPWR final_adder.U$$303/X sky130_fd_sc_hd__a21o_1
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$314 final_adder.U$$314/A final_adder.U$$314/B VGND VGND VPWR VPWR
+ final_adder.U$$348/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$325 final_adder.U$$324/A final_adder.U$$265/X final_adder.U$$267/X
+ VGND VGND VPWR VPWR final_adder.U$$325/X sky130_fd_sc_hd__a21o_1
Xrepeater540 U$$2733/A2 VGND VGND VPWR VPWR U$$2729/A2 sky130_fd_sc_hd__buf_4
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$336 final_adder.U$$336/A final_adder.U$$336/B VGND VGND VPWR VPWR
+ final_adder.U$$360/B sky130_fd_sc_hd__and2_2
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$347 final_adder.U$$346/A final_adder.U$$309/X final_adder.U$$311/X
+ VGND VGND VPWR VPWR ANTENNA_10/DIODE sky130_fd_sc_hd__a21o_1
Xrepeater551 U$$2437/A2 VGND VGND VPWR VPWR U$$2435/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$358 final_adder.U$$358/A final_adder.U$$358/B VGND VGND VPWR VPWR
+ final_adder.U$$370/A sky130_fd_sc_hd__and2_1
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater562 U$$2302/A2 VGND VGND VPWR VPWR U$$2298/A2 sky130_fd_sc_hd__buf_6
XU$$208 U$$208/A U$$216/B VGND VGND VPWR VPWR U$$208/X sky130_fd_sc_hd__xor2_1
Xrepeater573 U$$2185/A2 VGND VGND VPWR VPWR U$$2189/A2 sky130_fd_sc_hd__buf_6
XFILLER_38_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$369 final_adder.U$$354/X final_adder.U$$638/B final_adder.U$$355/X
+ VGND VGND VPWR VPWR final_adder.U$$654/B sky130_fd_sc_hd__a21o_4
Xrepeater584 U$$1851/A2 VGND VGND VPWR VPWR U$$1843/A2 sky130_fd_sc_hd__buf_6
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$219 U$$493/A1 U$$219/A2 U$$358/A1 U$$219/B2 VGND VGND VPWR VPWR U$$220/A sky130_fd_sc_hd__a22o_1
XFILLER_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater595 U$$1768/A2 VGND VGND VPWR VPWR U$$1762/A2 sky130_fd_sc_hd__buf_6
XFILLER_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_64_clk _535_/CLK VGND VGND VPWR VPWR _559_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_803 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2609_1737 VGND VGND VPWR VPWR U$$2609_1737/HI U$$2609/A1 sky130_fd_sc_hd__conb_1
XFILLER_129_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1108 U$$1370/A VGND VGND VPWR VPWR U$$1332/B sky130_fd_sc_hd__buf_6
XFILLER_119_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_111_1 U$$3687/X U$$3820/X U$$3953/X VGND VGND VPWR VPWR dadda_fa_4_112_1/B
+ dadda_fa_4_111_2/B sky130_fd_sc_hd__fa_1
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1119 _633_/Q VGND VGND VPWR VPWR U$$1203/B sky130_fd_sc_hd__clkbuf_8
XFILLER_181_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_104_0 U$$3806/X U$$3939/X U$$4072/X VGND VGND VPWR VPWR dadda_fa_4_105_0/B
+ dadda_fa_4_104_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_52_3 dadda_fa_3_52_3/A dadda_fa_3_52_3/B dadda_fa_3_52_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_1/B dadda_fa_4_52_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_209_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_68_3 U$$1473/X U$$1606/X U$$1739/X VGND VGND VPWR VPWR dadda_fa_1_69_6/CIN
+ dadda_fa_1_68_8/B sky130_fd_sc_hd__fa_1
XTAP_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_45_2 dadda_fa_3_45_2/A dadda_fa_3_45_2/B dadda_fa_3_45_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_1/A dadda_fa_4_45_2/B sky130_fd_sc_hd__fa_1
XFILLER_75_243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_38_1 dadda_fa_3_38_1/A dadda_fa_3_38_1/B dadda_fa_3_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_0/CIN dadda_fa_4_38_2/A sky130_fd_sc_hd__fa_1
XU$$720 U$$720/A U$$760/B VGND VGND VPWR VPWR U$$720/X sky130_fd_sc_hd__xor2_1
X_665_ _674_/CLK _665_/D VGND VGND VPWR VPWR _665_/Q sky130_fd_sc_hd__dfxtp_4
XU$$731 U$$731/A1 U$$759/A2 U$$733/A1 U$$759/B2 VGND VGND VPWR VPWR U$$732/A sky130_fd_sc_hd__a22o_1
XFILLER_91_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$742 U$$742/A U$$748/B VGND VGND VPWR VPWR U$$742/X sky130_fd_sc_hd__xor2_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_55_clk _535_/CLK VGND VGND VPWR VPWR _615_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_6_15_0 dadda_fa_6_15_0/A dadda_fa_6_15_0/B dadda_fa_6_15_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_16_0/B dadda_fa_7_15_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_189_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$753 U$$66/B1 U$$795/A2 U$$890/B1 U$$795/B2 VGND VGND VPWR VPWR U$$754/A sky130_fd_sc_hd__a22o_1
XFILLER_1_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$764 U$$764/A U$$766/B VGND VGND VPWR VPWR U$$764/X sky130_fd_sc_hd__xor2_1
X_596_ _596_/CLK _596_/D VGND VGND VPWR VPWR _596_/Q sky130_fd_sc_hd__dfxtp_4
XU$$775 U$$912/A1 U$$783/A2 U$$912/B1 U$$783/B2 VGND VGND VPWR VPWR U$$776/A sky130_fd_sc_hd__a22o_1
XFILLER_204_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$786 U$$786/A U$$821/A VGND VGND VPWR VPWR U$$786/X sky130_fd_sc_hd__xor2_1
XU$$797 U$$934/A1 U$$689/X U$$936/A1 U$$690/X VGND VGND VPWR VPWR U$$798/A sky130_fd_sc_hd__a22o_1
XFILLER_32_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_3_110_3 U$$4350/X U$$4483/X VGND VGND VPWR VPWR dadda_fa_4_111_1/CIN dadda_ha_3_110_3/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_204_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_532 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_3 _456_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_2_97_5 U$$4324/X U$$4457/X input253/X VGND VGND VPWR VPWR dadda_fa_3_98_2/A
+ dadda_fa_4_97_0/A sky130_fd_sc_hd__fa_2
Xrepeater1620 U$$4273/B1 VGND VGND VPWR VPWR U$$848/B1 sky130_fd_sc_hd__buf_6
XFILLER_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1631 U$$3451/A1 VGND VGND VPWR VPWR U$$985/A1 sky130_fd_sc_hd__buf_4
XFILLER_193_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1642 U$$3447/B1 VGND VGND VPWR VPWR U$$3584/B1 sky130_fd_sc_hd__buf_4
Xrepeater1653 _559_/Q VGND VGND VPWR VPWR U$$4404/B1 sky130_fd_sc_hd__buf_6
XFILLER_99_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1664 U$$2756/B1 VGND VGND VPWR VPWR U$$840/A1 sky130_fd_sc_hd__buf_6
XFILLER_67_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1675 U$$4400/A1 VGND VGND VPWR VPWR U$$2756/A1 sky130_fd_sc_hd__buf_8
XFILLER_140_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1686 _555_/Q VGND VGND VPWR VPWR U$$4259/B1 sky130_fd_sc_hd__buf_6
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1697 U$$3022/B1 VGND VGND VPWR VPWR U$$969/A1 sky130_fd_sc_hd__buf_4
XFILLER_112_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_40_1 U$$1949/X U$$2082/X U$$2215/X VGND VGND VPWR VPWR dadda_fa_3_41_0/CIN
+ dadda_fa_3_40_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_clk _369_/CLK VGND VGND VPWR VPWR _507_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_2_33_0 U$$73/X U$$206/X U$$339/X VGND VGND VPWR VPWR dadda_fa_3_34_0/B dadda_fa_3_33_2/B
+ sky130_fd_sc_hd__fa_1
XFILLER_19_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2160 U$$2160/A U$$2191/A VGND VGND VPWR VPWR U$$2160/X sky130_fd_sc_hd__xor2_1
XFILLER_74_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2171 U$$2171/A1 U$$2059/X U$$940/A1 U$$2060/X VGND VGND VPWR VPWR U$$2172/A sky130_fd_sc_hd__a22o_1
XU$$2182 U$$2182/A U$$2186/B VGND VGND VPWR VPWR U$$2182/X sky130_fd_sc_hd__xor2_1
XFILLER_168_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2193 _648_/Q VGND VGND VPWR VPWR U$$2195/B sky130_fd_sc_hd__inv_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1470 U$$2838/B1 U$$1474/A2 U$$2705/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1471/A
+ sky130_fd_sc_hd__a22o_1
XU$$1481 U$$1481/A U$$1487/B VGND VGND VPWR VPWR U$$1481/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1492 U$$2725/A1 U$$1500/A2 U$$2588/B1 U$$1500/B2 VGND VGND VPWR VPWR U$$1493/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_86_5 U$$3504/X U$$3637/X VGND VGND VPWR VPWR dadda_fa_2_87_4/B dadda_fa_3_86_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_163_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_3 U$$2704/X U$$2837/X U$$2970/X VGND VGND VPWR VPWR dadda_fa_2_86_3/B
+ dadda_fa_2_85_5/B sky130_fd_sc_hd__fa_1
XFILLER_131_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_62_2 dadda_fa_4_62_2/A dadda_fa_4_62_2/B dadda_fa_4_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/CIN dadda_fa_5_62_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_78_2 U$$2025/X U$$2158/X U$$2291/X VGND VGND VPWR VPWR dadda_fa_2_79_1/A
+ dadda_fa_2_78_4/A sky130_fd_sc_hd__fa_1
XFILLER_106_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_55_1 dadda_fa_4_55_1/A dadda_fa_4_55_1/B dadda_fa_4_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/B dadda_fa_5_55_1/B sky130_fd_sc_hd__fa_1
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$100 _524_/Q _396_/Q VGND VGND VPWR VPWR final_adder.U$$595/B1 final_adder.U$$722/A
+ sky130_fd_sc_hd__ha_1
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_32_0 dadda_fa_7_32_0/A dadda_fa_7_32_0/B dadda_fa_7_32_0/CIN VGND VGND
+ VPWR VPWR _457_/D _328_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$111 _535_/Q _407_/Q VGND VGND VPWR VPWR final_adder.U$$239/B1 final_adder.U$$733/A
+ sky130_fd_sc_hd__ha_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$122 _546_/Q _418_/Q VGND VGND VPWR VPWR final_adder.U$$617/B1 final_adder.U$$744/A
+ sky130_fd_sc_hd__ha_2
XFILLER_44_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_48_0 dadda_fa_4_48_0/A dadda_fa_4_48_0/B dadda_fa_4_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/A dadda_fa_5_48_1/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$133 final_adder.U$$627/A final_adder.U$$499/B1 final_adder.U$$5/COUT
+ VGND VGND VPWR VPWR final_adder.U$$133/X sky130_fd_sc_hd__a21o_1
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$144 final_adder.U$$639/A final_adder.U$$638/A VGND VGND VPWR VPWR
+ final_adder.U$$264/B sky130_fd_sc_hd__and2_1
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$155 final_adder.U$$649/A final_adder.U$$521/B1 final_adder.U$$155/B1
+ VGND VGND VPWR VPWR final_adder.U$$155/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$166 final_adder.U$$661/A final_adder.U$$660/A VGND VGND VPWR VPWR
+ final_adder.U$$274/A sky130_fd_sc_hd__and2_1
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$177 final_adder.U$$671/A final_adder.U$$543/B1 final_adder.U$$177/B1
+ VGND VGND VPWR VPWR final_adder.U$$177/X sky130_fd_sc_hd__a21o_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_991 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$188 final_adder.U$$683/A final_adder.U$$682/A VGND VGND VPWR VPWR
+ final_adder.U$$286/B sky130_fd_sc_hd__and2_1
XFILLER_166_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater392 U$$963/X VGND VGND VPWR VPWR U$$1065/A2 sky130_fd_sc_hd__buf_6
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$199 final_adder.U$$693/A final_adder.U$$565/B1 final_adder.U$$199/B1
+ VGND VGND VPWR VPWR final_adder.U$$199/X sky130_fd_sc_hd__a21o_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk _479_/CLK VGND VGND VPWR VPWR _234_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_450_ _451_/CLK _450_/D VGND VGND VPWR VPWR _450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_381_ _510_/CLK _381_/D VGND VGND VPWR VPWR _381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_73_1 U$$1084/X U$$1217/X U$$1350/X VGND VGND VPWR VPWR dadda_fa_1_74_7/CIN
+ dadda_fa_1_73_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_209_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_50_0 dadda_fa_3_50_0/A dadda_fa_3_50_0/B dadda_fa_3_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_0/B dadda_fa_4_50_1/CIN sky130_fd_sc_hd__fa_1
Xinput140 c[10] VGND VGND VPWR VPWR input140/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_0_66_0 _617_/Q U$$272/X U$$405/X VGND VGND VPWR VPWR dadda_fa_1_67_5/B dadda_fa_1_66_7/B
+ sky130_fd_sc_hd__fa_1
Xinput151 c[11] VGND VGND VPWR VPWR input151/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput162 c[14] VGND VGND VPWR VPWR input162/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput173 c[24] VGND VGND VPWR VPWR input173/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4447_1802 VGND VGND VPWR VPWR U$$4447_1802/HI U$$4447/B sky130_fd_sc_hd__conb_1
Xinput184 c[34] VGND VGND VPWR VPWR input184/X sky130_fd_sc_hd__clkbuf_4
XTAP_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput195 c[44] VGND VGND VPWR VPWR input195/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_28_clk _432_/CLK VGND VGND VPWR VPWR _213_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$550 U$$685/A VGND VGND VPWR VPWR U$$550/Y sky130_fd_sc_hd__inv_1
XFILLER_189_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_972 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_648_ _648_/CLK _648_/D VGND VGND VPWR VPWR _648_/Q sky130_fd_sc_hd__dfxtp_1
XU$$561 U$$561/A U$$589/B VGND VGND VPWR VPWR U$$561/X sky130_fd_sc_hd__xor2_1
XFILLER_205_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$572 U$$22/B1 U$$574/A2 U$$26/A1 U$$574/B2 VGND VGND VPWR VPWR U$$573/A sky130_fd_sc_hd__a22o_1
XFILLER_205_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$583 U$$583/A U$$659/B VGND VGND VPWR VPWR U$$583/X sky130_fd_sc_hd__xor2_1
XU$$594 U$$729/B1 U$$622/A2 U$$596/A1 U$$622/B2 VGND VGND VPWR VPWR U$$595/A sky130_fd_sc_hd__a22o_1
XFILLER_44_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_579_ _582_/CLK _579_/D VGND VGND VPWR VPWR _579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1069 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_362 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_95_2 U$$3389/X U$$3522/X U$$3655/X VGND VGND VPWR VPWR dadda_fa_3_96_1/A
+ dadda_fa_3_95_3/A sky130_fd_sc_hd__fa_1
XFILLER_172_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1450 _584_/Q VGND VGND VPWR VPWR U$$4045/A1 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_5_72_1 dadda_fa_5_72_1/A dadda_fa_5_72_1/B dadda_fa_5_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_73_0/B dadda_fa_7_72_0/A sky130_fd_sc_hd__fa_1
Xrepeater1461 U$$3493/A1 VGND VGND VPWR VPWR U$$66/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_88_1 U$$3907/X U$$4040/X U$$4173/X VGND VGND VPWR VPWR dadda_fa_3_89_0/CIN
+ dadda_fa_3_88_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_193_1050 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1472 U$$4176/A1 VGND VGND VPWR VPWR U$$3902/A1 sky130_fd_sc_hd__buf_4
XFILLER_113_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1483 U$$1843/A1 VGND VGND VPWR VPWR U$$882/B1 sky130_fd_sc_hd__buf_6
XFILLER_207_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1494 _578_/Q VGND VGND VPWR VPWR U$$3485/A1 sky130_fd_sc_hd__buf_6
XFILLER_28_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_65_0 dadda_fa_5_65_0/A dadda_fa_5_65_0/B dadda_fa_5_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_66_0/A dadda_fa_6_65_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_87 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_8 dadda_fa_1_64_8/A dadda_fa_1_64_8/B dadda_fa_1_64_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_3/A dadda_fa_3_64_0/A sky130_fd_sc_hd__fa_1
XFILLER_55_703 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_57_7 input209/X dadda_fa_1_57_7/B dadda_fa_1_57_7/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_58_2/CIN dadda_fa_2_57_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_4_0 U$$281/X U$$319/B input201/X VGND VGND VPWR VPWR dadda_fa_7_5_0/B
+ dadda_fa_7_4_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_90_1 U$$2182/X U$$2315/X U$$2448/X VGND VGND VPWR VPWR dadda_fa_2_91_4/B
+ dadda_fa_2_90_5/B sky130_fd_sc_hd__fa_1
XFILLER_2_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_83_0 U$$1369/Y U$$1503/X U$$1636/X VGND VGND VPWR VPWR dadda_fa_2_84_1/CIN
+ dadda_fa_2_83_4/A sky130_fd_sc_hd__fa_1
XFILLER_132_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4309 U$$4444/B1 U$$4335/A2 U$$4446/B1 U$$4311/B2 VGND VGND VPWR VPWR U$$4310/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3608 U$$4293/A1 U$$3612/A2 U$$4158/A1 U$$3612/B2 VGND VGND VPWR VPWR U$$3609/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3619 U$$3619/A U$$3627/B VGND VGND VPWR VPWR U$$3619/X sky130_fd_sc_hd__xor2_1
XFILLER_18_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_371 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2907 U$$3042/B1 U$$2959/A2 U$$2909/A1 U$$2959/B2 VGND VGND VPWR VPWR U$$2908/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2918 U$$2918/A U$$2944/B VGND VGND VPWR VPWR U$$2918/X sky130_fd_sc_hd__xor2_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_502_ _503_/CLK _502_/D VGND VGND VPWR VPWR _502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2929 U$$4436/A1 U$$2929/A2 U$$4436/B1 U$$2929/B2 VGND VGND VPWR VPWR U$$2930/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_212 _186_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 _187_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 _188_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_245 _194_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ _445_/CLK _433_/D VGND VGND VPWR VPWR _433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_278 _212_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_289 _214_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_364_ _494_/CLK _364_/D VGND VGND VPWR VPWR _364_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_295_ _615_/CLK _295_/D VGND VGND VPWR VPWR _295_/Q sky130_fd_sc_hd__dfxtp_1
XU$$4477_1817 VGND VGND VPWR VPWR U$$4477_1817/HI U$$4477/B sky130_fd_sc_hd__conb_1
XFILLER_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_82_0 dadda_fa_6_82_0/A dadda_fa_6_82_0/B dadda_fa_6_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_83_0/B dadda_fa_7_82_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_98_0 input254/X dadda_fa_3_98_0/B dadda_fa_3_98_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_99_0/B dadda_fa_4_98_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_155_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_674 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_364 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$380 U$$515/B1 U$$384/A2 U$$517/B1 U$$384/B2 VGND VGND VPWR VPWR U$$381/A sky130_fd_sc_hd__a22o_1
XFILLER_205_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$391 U$$391/A U$$393/B VGND VGND VPWR VPWR U$$391/X sky130_fd_sc_hd__xor2_1
XFILLER_178_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_clk _442_/CLK VGND VGND VPWR VPWR _445_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1280 U$$3539/A1 VGND VGND VPWR VPWR U$$2717/A1 sky130_fd_sc_hd__buf_6
Xrepeater1291 U$$3124/A1 VGND VGND VPWR VPWR U$$382/B1 sky130_fd_sc_hd__buf_8
XFILLER_102_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_5 U$$4298/B input215/X dadda_fa_1_62_5/CIN VGND VGND VPWR VPWR dadda_fa_2_63_2/A
+ dadda_fa_2_62_5/A sky130_fd_sc_hd__fa_1
XFILLER_80_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_55_4 U$$2378/X U$$2511/X U$$2644/X VGND VGND VPWR VPWR dadda_fa_2_56_1/CIN
+ dadda_fa_2_55_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_48_3 U$$1300/X U$$1433/X U$$1566/X VGND VGND VPWR VPWR dadda_fa_2_49_2/A
+ dadda_fa_2_48_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_43_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_25_2 dadda_fa_4_25_2/A dadda_fa_4_25_2/B dadda_fa_4_25_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/CIN dadda_fa_5_25_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_18_1 input166/X dadda_fa_4_18_1/B dadda_fa_4_18_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_5_19_0/B dadda_fa_5_18_1/B sky130_fd_sc_hd__fa_2
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_693 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4106 U$$4106/A U$$4109/A VGND VGND VPWR VPWR U$$4106/X sky130_fd_sc_hd__xor2_1
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_3_21_3 U$$1246/X U$$1379/X VGND VGND VPWR VPWR dadda_fa_4_22_1/B dadda_ha_3_21_3/SUM
+ sky130_fd_sc_hd__ha_1
XU$$4117 U$$4117/A U$$4141/B VGND VGND VPWR VPWR U$$4117/X sky130_fd_sc_hd__xor2_1
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4128 U$$4402/A1 U$$4226/A2 _558_/Q U$$4226/B2 VGND VGND VPWR VPWR U$$4129/A sky130_fd_sc_hd__a22o_1
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4139 U$$4139/A U$$4175/B VGND VGND VPWR VPWR U$$4139/X sky130_fd_sc_hd__xor2_1
XFILLER_59_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3405 U$$3405/A U$$3407/B VGND VGND VPWR VPWR U$$3405/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3416 U$$3551/B1 U$$3292/X U$$4514/A1 U$$3293/X VGND VGND VPWR VPWR U$$3417/A sky130_fd_sc_hd__a22o_1
XFILLER_46_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3427 _667_/Q VGND VGND VPWR VPWR U$$3427/Y sky130_fd_sc_hd__inv_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3438 U$$3438/A U$$3490/B VGND VGND VPWR VPWR U$$3438/X sky130_fd_sc_hd__xor2_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2704 U$$2704/A U$$2706/B VGND VGND VPWR VPWR U$$2704/X sky130_fd_sc_hd__xor2_1
XU$$3449 U$$3584/B1 U$$3497/A2 U$$3451/A1 U$$3497/B2 VGND VGND VPWR VPWR U$$3450/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2715 U$$2715/A1 U$$2733/A2 U$$2717/A1 U$$2733/B2 VGND VGND VPWR VPWR U$$2716/A
+ sky130_fd_sc_hd__a22o_1
XU$$2726 U$$2726/A U$$2730/B VGND VGND VPWR VPWR U$$2726/X sky130_fd_sc_hd__xor2_1
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2737 U$$2872/B1 U$$2607/X U$$2737/B1 U$$2608/X VGND VGND VPWR VPWR U$$2738/A sky130_fd_sc_hd__a22o_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2748 U$$3157/B1 U$$2798/A2 U$$3022/B1 U$$2798/B2 VGND VGND VPWR VPWR U$$2749/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_1 U$$446/X U$$579/X U$$712/X VGND VGND VPWR VPWR dadda_fa_4_21_0/CIN
+ dadda_fa_4_20_2/A sky130_fd_sc_hd__fa_1
XFILLER_15_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2759 U$$2759/A U$$2787/B VGND VGND VPWR VPWR U$$2759/X sky130_fd_sc_hd__xor2_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_416_ _547_/CLK _416_/D VGND VGND VPWR VPWR _416_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_347_ _475_/CLK _347_/D VGND VGND VPWR VPWR _347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_278_ _523_/CLK _278_/D VGND VGND VPWR VPWR _278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_527 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_700 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_72_4 dadda_fa_2_72_4/A dadda_fa_2_72_4/B dadda_fa_2_72_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/CIN dadda_fa_3_72_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_65_3 dadda_fa_2_65_3/A dadda_fa_2_65_3/B dadda_fa_2_65_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/B dadda_fa_3_65_3/B sky130_fd_sc_hd__fa_1
XFILLER_57_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater903 U$$4296/B VGND VGND VPWR VPWR U$$4298/B sky130_fd_sc_hd__buf_8
XFILLER_68_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater914 U$$4175/B VGND VGND VPWR VPWR U$$4141/B sky130_fd_sc_hd__buf_6
XFILLER_97_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater925 U$$4084/B VGND VGND VPWR VPWR U$$4109/A sky130_fd_sc_hd__buf_6
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater936 U$$3935/B VGND VGND VPWR VPWR U$$3917/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_58_2 dadda_fa_2_58_2/A dadda_fa_2_58_2/B dadda_fa_2_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/A dadda_fa_3_58_3/A sky130_fd_sc_hd__fa_1
XFILLER_37_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater947 _671_/Q VGND VGND VPWR VPWR U$$3836/A sky130_fd_sc_hd__buf_6
Xrepeater958 U$$3556/B VGND VGND VPWR VPWR U$$3506/B sky130_fd_sc_hd__buf_6
XFILLER_110_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_35_1 dadda_fa_5_35_1/A dadda_fa_5_35_1/B dadda_fa_5_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_36_0/B dadda_fa_7_35_0/A sky130_fd_sc_hd__fa_1
Xrepeater969 U$$3407/B VGND VGND VPWR VPWR U$$3363/B sky130_fd_sc_hd__buf_8
XFILLER_204_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_28_0 dadda_fa_5_28_0/A dadda_fa_5_28_0/B dadda_fa_5_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_29_0/A dadda_fa_6_28_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_209_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3950 U$$4087/A1 U$$3968/A2 U$$4087/B1 U$$3968/B2 VGND VGND VPWR VPWR U$$3951/A
+ sky130_fd_sc_hd__a22o_1
XU$$3961 U$$3961/A U$$3965/B VGND VGND VPWR VPWR U$$3961/X sky130_fd_sc_hd__xor2_1
XFILLER_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3972 U$$3973/A VGND VGND VPWR VPWR U$$3972/Y sky130_fd_sc_hd__inv_1
XFILLER_24_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3983 U$$4394/A1 U$$4005/A2 U$$4396/A1 U$$4005/B2 VGND VGND VPWR VPWR U$$3984/A
+ sky130_fd_sc_hd__a22o_1
XU$$3994 U$$3994/A U$$3994/B VGND VGND VPWR VPWR U$$3994/X sky130_fd_sc_hd__xor2_1
XFILLER_91_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_663 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_102_0 dadda_fa_5_102_0/A dadda_fa_5_102_0/B dadda_fa_5_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_103_0/A dadda_fa_6_102_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_482 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput263 _273_/Q VGND VGND VPWR VPWR o[105] sky130_fd_sc_hd__buf_2
XFILLER_173_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput274 _283_/Q VGND VGND VPWR VPWR o[115] sky130_fd_sc_hd__buf_2
XFILLER_160_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput285 _293_/Q VGND VGND VPWR VPWR o[125] sky130_fd_sc_hd__buf_2
XFILLER_142_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput296 _169_/Q VGND VGND VPWR VPWR o[1] sky130_fd_sc_hd__buf_2
XFILLER_59_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_60_2 U$$2787/X U$$2920/X U$$3053/X VGND VGND VPWR VPWR dadda_fa_2_61_1/A
+ dadda_fa_2_60_4/A sky130_fd_sc_hd__fa_1
XFILLER_75_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_53_1 U$$778/X U$$911/X U$$1044/X VGND VGND VPWR VPWR dadda_fa_2_54_0/CIN
+ dadda_fa_2_53_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_30_0 dadda_fa_4_30_0/A dadda_fa_4_30_0/B dadda_fa_4_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/A dadda_fa_5_30_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_46_0 U$$99/X U$$232/X U$$365/X VGND VGND VPWR VPWR dadda_fa_2_47_1/CIN
+ dadda_fa_2_46_4/A sky130_fd_sc_hd__fa_1
XFILLER_56_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_201_ _478_/CLK _201_/D VGND VGND VPWR VPWR _201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_438 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_82_3 dadda_fa_3_82_3/A dadda_fa_3_82_3/B dadda_fa_3_82_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_1/B dadda_fa_4_82_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_75_2 dadda_fa_3_75_2/A dadda_fa_3_75_2/B dadda_fa_3_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_1/A dadda_fa_4_75_2/B sky130_fd_sc_hd__fa_1
XFILLER_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_68_1 dadda_fa_3_68_1/A dadda_fa_3_68_1/B dadda_fa_3_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_0/CIN dadda_fa_4_68_2/A sky130_fd_sc_hd__fa_1
XFILLER_78_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_45_0 dadda_fa_6_45_0/A dadda_fa_6_45_0/B dadda_fa_6_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_46_0/B dadda_fa_7_45_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3202 U$$3202/A U$$3236/B VGND VGND VPWR VPWR U$$3202/X sky130_fd_sc_hd__xor2_1
XU$$3213 U$$3213/A1 U$$3215/A2 U$$3352/A1 U$$3215/B2 VGND VGND VPWR VPWR U$$3214/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3224 U$$3224/A U$$3232/B VGND VGND VPWR VPWR U$$3224/X sky130_fd_sc_hd__xor2_1
XU$$3235 U$$3372/A1 U$$3235/A2 U$$3374/A1 U$$3235/B2 VGND VGND VPWR VPWR U$$3236/A
+ sky130_fd_sc_hd__a22o_1
XU$$2501 U$$2501/A U$$2517/B VGND VGND VPWR VPWR U$$2501/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$17 _441_/Q _313_/Q VGND VGND VPWR VPWR final_adder.U$$145/B1 final_adder.U$$639/A
+ sky130_fd_sc_hd__ha_2
XFILLER_62_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$28 _452_/Q _324_/Q VGND VGND VPWR VPWR final_adder.U$$523/B1 final_adder.U$$650/A
+ sky130_fd_sc_hd__ha_2
XFILLER_111_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3246 U$$3246/A U$$3276/B VGND VGND VPWR VPWR U$$3246/X sky130_fd_sc_hd__xor2_1
XU$$3257 _601_/Q U$$3263/A2 _602_/Q U$$3263/B2 VGND VGND VPWR VPWR U$$3258/A sky130_fd_sc_hd__a22o_1
XU$$2512 U$$4154/B1 U$$2566/A2 U$$4156/B1 U$$2566/B2 VGND VGND VPWR VPWR U$$2513/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$39 _463_/Q _335_/Q VGND VGND VPWR VPWR final_adder.U$$167/B1 final_adder.U$$661/A
+ sky130_fd_sc_hd__ha_1
XU$$3268 U$$3268/A U$$3272/B VGND VGND VPWR VPWR U$$3268/X sky130_fd_sc_hd__xor2_1
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2523 U$$2523/A U$$2531/B VGND VGND VPWR VPWR U$$2523/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_104_2 dadda_fa_4_104_2/A dadda_fa_4_104_2/B dadda_fa_4_104_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/CIN dadda_fa_5_104_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2534 U$$3902/B1 U$$2470/X U$$3769/A1 U$$2471/X VGND VGND VPWR VPWR U$$2535/A sky130_fd_sc_hd__a22o_1
XU$$3279 U$$3551/B1 U$$3283/A2 U$$3281/A1 U$$3283/B2 VGND VGND VPWR VPWR U$$3280/A
+ sky130_fd_sc_hd__a22o_1
XU$$1800 U$$1800/A U$$1852/B VGND VGND VPWR VPWR U$$1800/X sky130_fd_sc_hd__xor2_1
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2545 U$$2545/A U$$2567/B VGND VGND VPWR VPWR U$$2545/X sky130_fd_sc_hd__xor2_1
XU$$2556 U$$3652/A1 U$$2588/A2 U$$914/A1 U$$2588/B2 VGND VGND VPWR VPWR U$$2557/A
+ sky130_fd_sc_hd__a22o_1
XU$$1811 U$$715/A1 U$$1851/A2 U$$715/B1 U$$1851/B2 VGND VGND VPWR VPWR U$$1812/A sky130_fd_sc_hd__a22o_1
XFILLER_34_558 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1822 U$$1822/A U$$1870/B VGND VGND VPWR VPWR U$$1822/X sky130_fd_sc_hd__xor2_1
XFILLER_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2567 U$$2567/A U$$2567/B VGND VGND VPWR VPWR U$$2567/X sky130_fd_sc_hd__xor2_1
XU$$1833 U$$52/A1 U$$1851/A2 U$$3342/A1 U$$1851/B2 VGND VGND VPWR VPWR U$$1834/A sky130_fd_sc_hd__a22o_1
XU$$2578 U$$3674/A1 U$$2580/A2 U$$2717/A1 U$$2580/B2 VGND VGND VPWR VPWR U$$2579/A
+ sky130_fd_sc_hd__a22o_1
XU$$1844 U$$1844/A U$$1844/B VGND VGND VPWR VPWR U$$1844/X sky130_fd_sc_hd__xor2_1
XU$$2589 U$$2589/A U$$2597/B VGND VGND VPWR VPWR U$$2589/X sky130_fd_sc_hd__xor2_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1855 U$$3362/A1 U$$1855/A2 U$$3362/B1 U$$1855/B2 VGND VGND VPWR VPWR U$$1856/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1866 U$$1866/A U$$1870/B VGND VGND VPWR VPWR U$$1866/X sky130_fd_sc_hd__xor2_1
XFILLER_159_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1877 U$$3245/B1 U$$1907/A2 U$$3112/A1 U$$1907/B2 VGND VGND VPWR VPWR U$$1878/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1888 U$$1888/A U$$1917/A VGND VGND VPWR VPWR U$$1888/X sky130_fd_sc_hd__xor2_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1899 U$$392/A1 U$$1909/A2 U$$3132/B1 U$$1909/B2 VGND VGND VPWR VPWR U$$1900/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_118_0 dadda_fa_7_118_0/A dadda_fa_7_118_0/B dadda_fa_7_118_0/CIN VGND
+ VGND VPWR VPWR _543_/D _414_/D sky130_fd_sc_hd__fa_1
XFILLER_119_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_786 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_70_1 dadda_fa_2_70_1/A dadda_fa_2_70_1/B dadda_fa_2_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_0/CIN dadda_fa_3_70_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_338 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_63_0 dadda_fa_2_63_0/A dadda_fa_2_63_0/B dadda_fa_2_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_0/B dadda_fa_3_63_2/B sky130_fd_sc_hd__fa_1
XFILLER_111_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater700 U$$4071/B2 VGND VGND VPWR VPWR U$$4065/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$507 final_adder.U$$634/A final_adder.U$$634/B final_adder.U$$507/B1
+ VGND VGND VPWR VPWR final_adder.U$$635/B sky130_fd_sc_hd__a21o_1
Xrepeater711 U$$3823/B2 VGND VGND VPWR VPWR U$$3769/B2 sky130_fd_sc_hd__buf_6
Xrepeater722 U$$3674/B2 VGND VGND VPWR VPWR U$$3688/B2 sky130_fd_sc_hd__buf_6
XFILLER_97_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$529 final_adder.U$$656/A final_adder.U$$656/B final_adder.U$$529/B1
+ VGND VGND VPWR VPWR final_adder.U$$657/B sky130_fd_sc_hd__a21o_1
Xrepeater733 U$$3430/X VGND VGND VPWR VPWR U$$3555/B2 sky130_fd_sc_hd__buf_6
Xrepeater744 U$$3231/B2 VGND VGND VPWR VPWR U$$3215/B2 sky130_fd_sc_hd__buf_4
XFILLER_96_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater755 U$$3132/B2 VGND VGND VPWR VPWR U$$3120/B2 sky130_fd_sc_hd__buf_6
Xrepeater766 U$$2882/X VGND VGND VPWR VPWR U$$2973/B2 sky130_fd_sc_hd__buf_6
Xrepeater777 U$$2798/B2 VGND VGND VPWR VPWR U$$2788/B2 sky130_fd_sc_hd__buf_4
Xrepeater788 U$$2733/B2 VGND VGND VPWR VPWR U$$2729/B2 sky130_fd_sc_hd__buf_4
XU$$4470 U$$4470/A1 U$$4388/X U$$4472/A1 U$$4480/B2 VGND VGND VPWR VPWR U$$4471/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater799 U$$2437/B2 VGND VGND VPWR VPWR U$$2435/B2 sky130_fd_sc_hd__buf_4
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4481 U$$4481/A U$$4481/B VGND VGND VPWR VPWR U$$4481/X sky130_fd_sc_hd__xor2_1
XU$$4492 U$$930/A1 U$$4388/X U$$932/A1 U$$4496/B2 VGND VGND VPWR VPWR U$$4493/A sky130_fd_sc_hd__a22o_1
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3780 U$$3780/A U$$3800/B VGND VGND VPWR VPWR U$$3780/X sky130_fd_sc_hd__xor2_1
XFILLER_92_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3791 _594_/Q U$$3795/A2 U$$3791/B1 U$$3795/B2 VGND VGND VPWR VPWR U$$3792/A sky130_fd_sc_hd__a22o_1
XFILLER_197_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_919 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_92_2 dadda_fa_4_92_2/A dadda_fa_4_92_2/B dadda_fa_4_92_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/CIN dadda_fa_5_92_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_146_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_85_1 dadda_fa_4_85_1/A dadda_fa_4_85_1/B dadda_fa_4_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/B dadda_fa_5_85_1/B sky130_fd_sc_hd__fa_1
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_62_0 dadda_fa_7_62_0/A dadda_fa_7_62_0/B dadda_fa_7_62_0/CIN VGND VGND
+ VPWR VPWR _487_/D _358_/D sky130_fd_sc_hd__fa_1
XFILLER_122_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_78_0 dadda_fa_4_78_0/A dadda_fa_4_78_0/B dadda_fa_4_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/A dadda_fa_5_78_1/A sky130_fd_sc_hd__fa_1
XFILLER_0_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$902 U$$80/A1 U$$906/A2 U$$80/B1 U$$906/B2 VGND VGND VPWR VPWR U$$903/A sky130_fd_sc_hd__a22o_1
XU$$913 U$$913/A U$$958/A VGND VGND VPWR VPWR U$$913/X sky130_fd_sc_hd__xor2_1
XU$$924 U$$924/A1 U$$924/A2 U$$924/B1 U$$924/B2 VGND VGND VPWR VPWR U$$925/A sky130_fd_sc_hd__a22o_1
XFILLER_84_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$935 U$$935/A U$$935/B VGND VGND VPWR VPWR U$$935/X sky130_fd_sc_hd__xor2_1
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$946 U$$946/A1 U$$948/A2 U$$946/B1 U$$948/B2 VGND VGND VPWR VPWR U$$947/A sky130_fd_sc_hd__a22o_1
XU$$957 U$$957/A U$$958/A VGND VGND VPWR VPWR U$$957/X sky130_fd_sc_hd__xor2_1
XU$$968 U$$968/A U$$994/B VGND VGND VPWR VPWR U$$968/X sky130_fd_sc_hd__xor2_1
XU$$1107 U$$1107/A U$$1151/B VGND VGND VPWR VPWR U$$1107/X sky130_fd_sc_hd__xor2_1
XFILLER_189_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$979 U$$20/A1 U$$979/A2 U$$20/B1 U$$979/B2 VGND VGND VPWR VPWR U$$980/A sky130_fd_sc_hd__a22o_1
XU$$1118 U$$22/A1 U$$1150/A2 U$$24/A1 U$$1150/B2 VGND VGND VPWR VPWR U$$1119/A sky130_fd_sc_hd__a22o_1
XU$$1129 U$$1129/A U$$1195/B VGND VGND VPWR VPWR U$$1129/X sky130_fd_sc_hd__xor2_1
XFILLER_203_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_80_0 dadda_fa_3_80_0/A dadda_fa_3_80_0/B dadda_fa_3_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_0/B dadda_fa_4_80_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_338 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3010 U$$3010/A _659_/Q VGND VGND VPWR VPWR U$$3010/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_42_5 dadda_fa_2_42_5/A dadda_fa_2_42_5/B dadda_fa_2_42_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_43_2/A dadda_fa_4_42_0/A sky130_fd_sc_hd__fa_2
XFILLER_47_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3021 U$$3021/A U$$3065/B VGND VGND VPWR VPWR U$$3021/X sky130_fd_sc_hd__xor2_1
XU$$3032 U$$3578/B1 U$$3046/A2 U$$3445/A1 U$$3046/B2 VGND VGND VPWR VPWR U$$3033/A
+ sky130_fd_sc_hd__a22o_1
XU$$3043 U$$3043/A U$$3083/B VGND VGND VPWR VPWR U$$3043/X sky130_fd_sc_hd__xor2_1
XFILLER_93_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3054 U$$3054/A1 U$$3054/A2 U$$3193/A1 U$$3054/B2 VGND VGND VPWR VPWR U$$3055/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_35_4 U$$1939/X U$$2072/X U$$2205/X VGND VGND VPWR VPWR dadda_fa_3_36_1/CIN
+ dadda_fa_3_35_3/CIN sky130_fd_sc_hd__fa_1
XU$$2320 _612_/Q U$$2326/A2 U$$2459/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2321/A sky130_fd_sc_hd__a22o_1
XU$$3065 U$$3065/A U$$3065/B VGND VGND VPWR VPWR U$$3065/X sky130_fd_sc_hd__xor2_1
XFILLER_35_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2331 U$$2466/A VGND VGND VPWR VPWR U$$2331/Y sky130_fd_sc_hd__inv_1
XU$$3076 U$$3896/B1 U$$3082/A2 U$$4448/A1 U$$3082/B2 VGND VGND VPWR VPWR U$$3077/A
+ sky130_fd_sc_hd__a22o_1
XU$$3087 U$$3087/A U$$3121/B VGND VGND VPWR VPWR U$$3087/X sky130_fd_sc_hd__xor2_1
XU$$2342 U$$2342/A U$$2366/B VGND VGND VPWR VPWR U$$2342/X sky130_fd_sc_hd__xor2_1
XU$$2353 U$$3584/B1 U$$2395/A2 U$$435/B1 U$$2395/B2 VGND VGND VPWR VPWR U$$2354/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3098 U$$3646/A1 U$$3110/A2 U$$4470/A1 U$$3110/B2 VGND VGND VPWR VPWR U$$3099/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2364 U$$2364/A U$$2388/B VGND VGND VPWR VPWR U$$2364/X sky130_fd_sc_hd__xor2_1
XU$$2375 U$$2375/A1 U$$2423/A2 U$$2375/B1 U$$2423/B2 VGND VGND VPWR VPWR U$$2376/A
+ sky130_fd_sc_hd__a22o_1
XU$$1630 U$$1630/A U$$1636/B VGND VGND VPWR VPWR U$$1630/X sky130_fd_sc_hd__xor2_1
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1641 U$$4105/B1 U$$1511/X U$$1641/B1 U$$1512/X VGND VGND VPWR VPWR U$$1642/A sky130_fd_sc_hd__a22o_1
XFILLER_61_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2386 U$$2386/A U$$2388/B VGND VGND VPWR VPWR U$$2386/X sky130_fd_sc_hd__xor2_1
XU$$2397 U$$3902/B1 U$$2437/A2 U$$3769/A1 U$$2437/B2 VGND VGND VPWR VPWR U$$2398/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1652 U$$2746/B1 U$$1684/A2 U$$695/A1 U$$1684/B2 VGND VGND VPWR VPWR U$$1653/A
+ sky130_fd_sc_hd__a22o_1
XU$$1663 U$$1663/A U$$1687/B VGND VGND VPWR VPWR U$$1663/X sky130_fd_sc_hd__xor2_1
XFILLER_50_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1674 U$$3042/B1 U$$1710/A2 U$$2909/A1 U$$1710/B2 VGND VGND VPWR VPWR U$$1675/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1685 U$$1685/A U$$1687/B VGND VGND VPWR VPWR U$$1685/X sky130_fd_sc_hd__xor2_1
XFILLER_203_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1696 U$$52/A1 U$$1740/A2 U$$52/B1 U$$1740/B2 VGND VGND VPWR VPWR U$$1697/A sky130_fd_sc_hd__a22o_1
XFILLER_124_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_95_0 dadda_fa_5_95_0/A dadda_fa_5_95_0/B dadda_fa_5_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_96_0/A dadda_fa_6_95_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_135_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_588 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$304 final_adder.U$$304/A final_adder.U$$304/B VGND VGND VPWR VPWR
+ final_adder.U$$344/B sky130_fd_sc_hd__and2_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$315 final_adder.U$$314/A final_adder.U$$245/X final_adder.U$$247/X
+ VGND VGND VPWR VPWR final_adder.U$$315/X sky130_fd_sc_hd__a21o_1
Xrepeater530 U$$2744/X VGND VGND VPWR VPWR U$$2798/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$326 final_adder.U$$326/A final_adder.U$$326/B VGND VGND VPWR VPWR
+ final_adder.U$$354/A sky130_fd_sc_hd__and2_1
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$337 final_adder.U$$336/A final_adder.U$$289/X final_adder.U$$291/X
+ VGND VGND VPWR VPWR final_adder.U$$337/X sky130_fd_sc_hd__a21o_2
Xrepeater541 U$$2607/X VGND VGND VPWR VPWR U$$2733/A2 sky130_fd_sc_hd__buf_4
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$348 final_adder.U$$348/A final_adder.U$$348/B VGND VGND VPWR VPWR
+ final_adder.U$$348/X sky130_fd_sc_hd__and2_1
Xrepeater552 U$$2387/A2 VGND VGND VPWR VPWR U$$2367/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$359 final_adder.U$$358/A final_adder.U$$333/X final_adder.U$$335/X
+ VGND VGND VPWR VPWR final_adder.U$$359/X sky130_fd_sc_hd__a21o_1
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater563 U$$2274/A2 VGND VGND VPWR VPWR U$$2302/A2 sky130_fd_sc_hd__buf_6
XU$$209 U$$72/A1 U$$217/A2 U$$74/A1 U$$217/B2 VGND VGND VPWR VPWR U$$210/A sky130_fd_sc_hd__a22o_1
Xrepeater574 U$$2059/X VGND VGND VPWR VPWR U$$2185/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater585 U$$1907/A2 VGND VGND VPWR VPWR U$$1851/A2 sky130_fd_sc_hd__buf_4
XFILLER_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater596 U$$1778/A2 VGND VGND VPWR VPWR U$$1768/A2 sky130_fd_sc_hd__buf_6
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_583 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1109 U$$1370/A VGND VGND VPWR VPWR U$$1369/A sky130_fd_sc_hd__buf_8
XFILLER_101_1031 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_931 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_111_2 U$$4086/X U$$4219/X U$$4352/X VGND VGND VPWR VPWR dadda_fa_4_112_1/CIN
+ dadda_fa_4_111_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_104_1 U$$4205/X U$$4338/X U$$4471/X VGND VGND VPWR VPWR dadda_fa_4_105_0/CIN
+ dadda_fa_4_104_2/A sky130_fd_sc_hd__fa_1
XFILLER_105_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_125_0 input157/X dadda_fa_6_125_0/B dadda_fa_6_125_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_126_0/B dadda_fa_7_125_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_68_4 U$$1872/X U$$2005/X U$$2138/X VGND VGND VPWR VPWR dadda_fa_1_69_7/A
+ dadda_fa_1_68_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_209_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_45_3 dadda_fa_3_45_3/A dadda_fa_3_45_3/B dadda_fa_3_45_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_1/B dadda_fa_4_45_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$710 U$$710/A U$$766/B VGND VGND VPWR VPWR U$$710/X sky130_fd_sc_hd__xor2_1
XTAP_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_38_2 dadda_fa_3_38_2/A dadda_fa_3_38_2/B dadda_fa_3_38_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_1/A dadda_fa_4_38_2/B sky130_fd_sc_hd__fa_1
X_664_ _674_/CLK _664_/D VGND VGND VPWR VPWR _664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$721 U$$856/B1 U$$759/A2 U$$997/A1 U$$759/B2 VGND VGND VPWR VPWR U$$722/A sky130_fd_sc_hd__a22o_1
XU$$732 U$$732/A U$$760/B VGND VGND VPWR VPWR U$$732/X sky130_fd_sc_hd__xor2_1
XU$$743 U$$880/A1 U$$747/A2 U$$745/A1 U$$747/B2 VGND VGND VPWR VPWR U$$744/A sky130_fd_sc_hd__a22o_1
XFILLER_204_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$754 U$$754/A U$$796/B VGND VGND VPWR VPWR U$$754/X sky130_fd_sc_hd__xor2_1
XFILLER_186_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$765 U$$900/B1 U$$765/A2 U$$82/A1 U$$765/B2 VGND VGND VPWR VPWR U$$766/A sky130_fd_sc_hd__a22o_1
X_595_ _596_/CLK _595_/D VGND VGND VPWR VPWR _595_/Q sky130_fd_sc_hd__dfxtp_4
XU$$776 U$$776/A U$$816/B VGND VGND VPWR VPWR U$$776/X sky130_fd_sc_hd__xor2_1
XFILLER_56_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$787 U$$924/A1 U$$809/A2 U$$924/B1 U$$809/B2 VGND VGND VPWR VPWR U$$788/A sky130_fd_sc_hd__a22o_1
XFILLER_95_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$798 U$$798/A U$$804/B VGND VGND VPWR VPWR U$$798/X sky130_fd_sc_hd__xor2_1
XFILLER_43_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1610 U$$4416/A1 VGND VGND VPWR VPWR U$$3181/B1 sky130_fd_sc_hd__buf_8
XANTENNA_4 _456_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1621 U$$987/A1 VGND VGND VPWR VPWR U$$28/A1 sky130_fd_sc_hd__buf_4
Xrepeater1632 U$$3312/B1 VGND VGND VPWR VPWR U$$3451/A1 sky130_fd_sc_hd__buf_6
Xrepeater1643 U$$3447/B1 VGND VGND VPWR VPWR U$$3175/A1 sky130_fd_sc_hd__buf_6
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1654 U$$20/A1 VGND VGND VPWR VPWR U$$2210/B1 sky130_fd_sc_hd__buf_6
Xrepeater1665 U$$2893/B1 VGND VGND VPWR VPWR U$$2756/B1 sky130_fd_sc_hd__buf_4
XFILLER_154_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1676 U$$3713/B1 VGND VGND VPWR VPWR U$$4400/A1 sky130_fd_sc_hd__buf_8
XFILLER_113_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3979_1759 VGND VGND VPWR VPWR U$$3979_1759/HI U$$3979/A1 sky130_fd_sc_hd__conb_1
Xrepeater1687 _554_/Q VGND VGND VPWR VPWR U$$4396/A1 sky130_fd_sc_hd__buf_8
XFILLER_99_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1698 U$$556/B1 VGND VGND VPWR VPWR U$$3022/B1 sky130_fd_sc_hd__buf_6
XFILLER_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_2_27_2 U$$859/X U$$992/X VGND VGND VPWR VPWR dadda_fa_3_28_2/CIN dadda_fa_4_27_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_94_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1059 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_40_2 U$$2348/X U$$2481/X U$$2614/X VGND VGND VPWR VPWR dadda_fa_3_41_1/A
+ dadda_fa_3_40_3/A sky130_fd_sc_hd__fa_1
XFILLER_94_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_33_1 U$$472/X U$$605/X U$$738/X VGND VGND VPWR VPWR dadda_fa_3_34_0/CIN
+ dadda_fa_3_33_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2150 U$$2150/A U$$2170/B VGND VGND VPWR VPWR U$$2150/X sky130_fd_sc_hd__xor2_1
XFILLER_34_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_10_0 U$$692/X U$$760/B input140/X VGND VGND VPWR VPWR dadda_fa_6_11_0/A
+ dadda_fa_6_10_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_179_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_26_0 U$$59/X U$$192/X U$$325/X VGND VGND VPWR VPWR dadda_fa_3_27_2/B dadda_fa_3_26_3/B
+ sky130_fd_sc_hd__fa_1
XU$$2161 U$$3255/B1 U$$2169/A2 U$$3122/A1 U$$2169/B2 VGND VGND VPWR VPWR U$$2162/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2172 U$$2172/A U$$2174/B VGND VGND VPWR VPWR U$$2172/X sky130_fd_sc_hd__xor2_1
XU$$2183 U$$2318/B1 U$$2185/A2 U$$3418/A1 U$$2185/B2 VGND VGND VPWR VPWR U$$2184/A
+ sky130_fd_sc_hd__a22o_1
XU$$2194 _649_/Q VGND VGND VPWR VPWR U$$2194/Y sky130_fd_sc_hd__inv_1
XU$$1460 U$$90/A1 U$$1474/A2 U$$92/A1 U$$1474/B2 VGND VGND VPWR VPWR U$$1461/A sky130_fd_sc_hd__a22o_1
XFILLER_50_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1471 U$$1471/A U$$1475/B VGND VGND VPWR VPWR U$$1471/X sky130_fd_sc_hd__xor2_1
XU$$1482 U$$2715/A1 U$$1500/A2 U$$525/A1 U$$1500/B2 VGND VGND VPWR VPWR U$$1483/A
+ sky130_fd_sc_hd__a22o_1
XU$$1493 U$$1493/A U$$1501/B VGND VGND VPWR VPWR U$$1493/X sky130_fd_sc_hd__xor2_1
XFILLER_124_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_85_4 U$$3103/X U$$3236/X U$$3369/X VGND VGND VPWR VPWR dadda_fa_2_86_3/CIN
+ dadda_fa_2_85_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_78_3 U$$2424/X U$$2557/X U$$2690/X VGND VGND VPWR VPWR dadda_fa_2_79_1/B
+ dadda_fa_2_78_4/B sky130_fd_sc_hd__fa_1
XFILLER_132_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_55_2 dadda_fa_4_55_2/A dadda_fa_4_55_2/B dadda_fa_4_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/CIN dadda_fa_5_55_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$101 _525_/Q _397_/Q VGND VGND VPWR VPWR final_adder.U$$229/B1 final_adder.U$$723/A
+ sky130_fd_sc_hd__ha_1
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$112 _536_/Q _408_/Q VGND VGND VPWR VPWR final_adder.U$$607/B1 ANTENNA_9/DIODE
+ sky130_fd_sc_hd__ha_4
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$123 _547_/Q _419_/Q VGND VGND VPWR VPWR final_adder.U$$251/B1 final_adder.U$$745/A
+ sky130_fd_sc_hd__ha_2
Xdadda_fa_4_48_1 dadda_fa_4_48_1/A dadda_fa_4_48_1/B dadda_fa_4_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/B dadda_fa_5_48_1/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$134 final_adder.U$$7/SUM final_adder.U$$628/A VGND VGND VPWR VPWR
+ final_adder.U$$258/A sky130_fd_sc_hd__and2_1
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$145 final_adder.U$$639/A final_adder.U$$511/B1 final_adder.U$$145/B1
+ VGND VGND VPWR VPWR final_adder.U$$145/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_7_25_0 dadda_fa_7_25_0/A dadda_fa_7_25_0/B dadda_fa_7_25_0/CIN VGND VGND
+ VPWR VPWR _450_/D _321_/D sky130_fd_sc_hd__fa_1
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$156 final_adder.U$$651/A final_adder.U$$650/A VGND VGND VPWR VPWR
+ final_adder.U$$270/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$167 final_adder.U$$661/A final_adder.U$$533/B1 final_adder.U$$167/B1
+ VGND VGND VPWR VPWR final_adder.U$$167/X sky130_fd_sc_hd__a21o_1
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$178 final_adder.U$$673/A final_adder.U$$672/A VGND VGND VPWR VPWR
+ final_adder.U$$280/A sky130_fd_sc_hd__and2_1
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$189 final_adder.U$$683/A final_adder.U$$555/B1 final_adder.U$$189/B1
+ VGND VGND VPWR VPWR final_adder.U$$189/X sky130_fd_sc_hd__a21o_1
Xrepeater393 U$$928/A2 VGND VGND VPWR VPWR U$$860/A2 sky130_fd_sc_hd__buf_4
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_380_ _510_/CLK _380_/D VGND VGND VPWR VPWR _380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_73_2 U$$1483/X U$$1616/X U$$1749/X VGND VGND VPWR VPWR dadda_fa_1_74_8/A
+ dadda_fa_2_73_0/A sky130_fd_sc_hd__fa_2
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput130 c[100] VGND VGND VPWR VPWR input130/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_691 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_50_1 dadda_fa_3_50_1/A dadda_fa_3_50_1/B dadda_fa_3_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_0/CIN dadda_fa_4_50_2/A sky130_fd_sc_hd__fa_1
XFILLER_0_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput141 c[110] VGND VGND VPWR VPWR input141/X sky130_fd_sc_hd__dlymetal6s2s_1
Xdadda_fa_0_66_1 U$$538/X U$$671/X U$$804/X VGND VGND VPWR VPWR dadda_fa_1_67_5/CIN
+ dadda_fa_1_66_7/CIN sky130_fd_sc_hd__fa_1
Xinput152 c[120] VGND VGND VPWR VPWR input152/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput163 c[15] VGND VGND VPWR VPWR input163/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput174 c[25] VGND VGND VPWR VPWR input174/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_3_43_0 dadda_fa_3_43_0/A dadda_fa_3_43_0/B dadda_fa_3_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_0/B dadda_fa_4_43_1/CIN sky130_fd_sc_hd__fa_1
Xinput185 c[35] VGND VGND VPWR VPWR input185/X sky130_fd_sc_hd__buf_4
XFILLER_76_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput196 c[45] VGND VGND VPWR VPWR input196/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_0_59_0 U$$125/X U$$258/X U$$391/X VGND VGND VPWR VPWR dadda_fa_1_60_6/B
+ dadda_fa_1_59_8/A sky130_fd_sc_hd__fa_1
XTAP_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$690 final_adder.U$$690/A final_adder.U$$690/B VGND VGND VPWR VPWR
+ _236_/D sky130_fd_sc_hd__xor2_4
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$540 U$$540/A _623_/Q VGND VGND VPWR VPWR U$$540/X sky130_fd_sc_hd__xor2_1
XFILLER_45_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_647_ _660_/CLK _647_/D VGND VGND VPWR VPWR _647_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$551 U$$685/A U$$551/B VGND VGND VPWR VPWR U$$551/X sky130_fd_sc_hd__and2_1
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$562 U$$562/A1 U$$574/A2 U$$973/B1 U$$574/B2 VGND VGND VPWR VPWR U$$563/A sky130_fd_sc_hd__a22o_1
XFILLER_189_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$573 U$$573/A U$$589/B VGND VGND VPWR VPWR U$$573/X sky130_fd_sc_hd__xor2_1
XFILLER_45_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$584 U$$719/B1 U$$600/A2 U$$584/B1 U$$600/B2 VGND VGND VPWR VPWR U$$585/A sky130_fd_sc_hd__a22o_1
XFILLER_189_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_578_ _582_/CLK _578_/D VGND VGND VPWR VPWR _578_/Q sky130_fd_sc_hd__dfxtp_4
XU$$595 U$$595/A U$$665/B VGND VGND VPWR VPWR U$$595/X sky130_fd_sc_hd__xor2_1
XFILLER_32_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_1097 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_971 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_100_0 dadda_fa_7_100_0/A dadda_fa_7_100_0/B dadda_fa_7_100_0/CIN VGND
+ VGND VPWR VPWR _525_/D _396_/D sky130_fd_sc_hd__fa_1
XFILLER_157_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_95_3 U$$3788/X U$$3921/X U$$4054/X VGND VGND VPWR VPWR dadda_fa_3_96_1/B
+ dadda_fa_3_95_3/B sky130_fd_sc_hd__fa_1
XFILLER_172_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1440 _585_/Q VGND VGND VPWR VPWR U$$4184/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_99_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1451 U$$3221/A1 VGND VGND VPWR VPWR U$$344/A1 sky130_fd_sc_hd__buf_4
XFILLER_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1462 U$$4450/B1 VGND VGND VPWR VPWR U$$3493/A1 sky130_fd_sc_hd__buf_6
XFILLER_154_1002 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_88_2 U$$4306/X U$$4439/X input243/X VGND VGND VPWR VPWR dadda_fa_3_89_1/A
+ dadda_fa_3_88_3/A sky130_fd_sc_hd__fa_1
Xrepeater1473 U$$4450/A1 VGND VGND VPWR VPWR U$$4176/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_207_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1484 U$$3213/A1 VGND VGND VPWR VPWR U$$1843/A1 sky130_fd_sc_hd__buf_4
XFILLER_67_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_65_1 dadda_fa_5_65_1/A dadda_fa_5_65_1/B dadda_fa_5_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_66_0/B dadda_fa_7_65_0/A sky130_fd_sc_hd__fa_1
Xrepeater1495 U$$334/A1 VGND VGND VPWR VPWR U$$60/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_58_0 dadda_fa_5_58_0/A dadda_fa_5_58_0/B dadda_fa_5_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_59_0/A dadda_fa_6_58_0/CIN sky130_fd_sc_hd__fa_2
.ends

