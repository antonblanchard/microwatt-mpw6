VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 14.090 2934.450 17.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 194.090 2934.450 197.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 374.090 2934.450 377.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 554.090 2934.450 557.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 734.090 2934.450 737.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 914.090 2934.450 917.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1094.090 2934.450 1097.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1274.090 2934.450 1277.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1454.090 2934.450 1457.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1634.090 2934.450 1637.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1814.090 2934.450 1817.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1994.090 2934.450 1997.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2174.090 2934.450 2177.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2354.090 2934.450 2357.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2534.090 2934.450 2537.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2714.090 2934.450 2717.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2894.090 2934.450 2897.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3074.090 2934.450 3077.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3254.090 2934.450 3257.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3434.090 2934.450 3437.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -9.470 12.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 -9.470 192.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 -9.470 372.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 -9.470 552.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 -9.470 732.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 -9.470 912.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 -9.470 1092.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 -9.470 1812.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 -9.470 1992.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 -9.470 2172.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 -9.470 2352.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 -9.470 2532.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 -9.470 2712.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2888.970 -9.470 2892.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 236.000 12.070 517.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 236.000 192.070 517.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 236.000 372.070 517.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 236.000 552.070 517.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 236.000 1812.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 236.000 1992.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 236.000 2172.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 236.000 2352.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 236.000 2532.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 236.000 2712.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2888.970 236.000 2892.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 1137.440 12.070 1584.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 1137.440 192.070 1584.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1137.440 372.070 1584.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 1137.440 552.070 1584.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 236.000 732.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 236.000 912.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 236.000 1092.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 -9.470 1272.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 -9.470 1452.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 -9.470 1632.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 1945.840 1812.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 1945.840 1992.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1945.840 2172.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 2203.680 12.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 2203.680 192.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2203.680 372.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2203.680 552.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 3488.640 732.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 3488.640 912.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 3488.640 1092.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 3488.640 1272.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 3488.640 1452.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 3488.640 1632.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 3488.640 1812.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 3488.640 1992.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 3488.640 2172.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 1945.840 2352.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 1945.840 2532.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 1945.840 2712.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2888.970 1945.840 2892.070 3529.150 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 32.930 2944.050 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 212.930 2944.050 216.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 392.930 2944.050 396.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 572.930 2944.050 576.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 752.930 2944.050 756.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 932.930 2944.050 936.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1112.930 2944.050 1116.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1292.930 2944.050 1296.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1472.930 2944.050 1476.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1652.930 2944.050 1656.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1832.930 2944.050 1836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2012.930 2944.050 2016.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2192.930 2944.050 2196.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2372.930 2944.050 2376.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2552.930 2944.050 2556.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2732.930 2944.050 2736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2912.930 2944.050 2916.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3092.930 2944.050 3096.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3272.930 2944.050 3276.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3452.930 2944.050 3456.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -19.070 30.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 -19.070 210.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 -19.070 390.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 -19.070 570.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 -19.070 750.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 -19.070 930.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 -19.070 1110.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 -19.070 1830.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 -19.070 2010.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 -19.070 2190.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 -19.070 2370.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 -19.070 2550.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 -19.070 2730.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.570 -19.070 2910.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 236.240 30.670 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 236.240 210.670 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 236.240 390.670 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 236.240 570.670 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 236.240 1830.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 236.240 2010.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 236.240 2190.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 236.240 2370.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 236.240 2550.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 236.240 2730.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.570 236.240 2910.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 1137.680 30.670 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 1137.680 210.670 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 1137.680 390.670 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 1137.680 570.670 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 236.240 750.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 236.240 930.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 236.240 1110.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 -19.070 1290.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 -19.070 1470.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 -19.070 1650.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 1946.080 1830.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 1946.080 2010.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 1946.080 2190.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 2203.920 30.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 2203.920 210.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 2203.920 390.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 2203.920 570.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 3488.880 750.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 3488.880 930.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 3488.880 1110.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 3488.880 1290.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 3488.880 1470.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 3488.880 1650.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 3488.880 1830.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 3488.880 2010.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 3488.880 2190.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 1946.080 2370.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 1946.080 2550.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 1946.080 2730.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.570 1946.080 2910.670 3538.750 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 51.530 2953.650 54.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 231.530 2953.650 234.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 411.530 2953.650 414.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 591.530 2953.650 594.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 771.530 2953.650 774.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 951.530 2953.650 954.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1131.530 2953.650 1134.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1311.530 2953.650 1314.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1491.530 2953.650 1494.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1671.530 2953.650 1674.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1851.530 2953.650 1854.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2031.530 2953.650 2034.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2211.530 2953.650 2214.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2391.530 2953.650 2394.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2571.530 2953.650 2574.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2751.530 2953.650 2754.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2931.530 2953.650 2934.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3111.530 2953.650 3114.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3291.530 2953.650 3294.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3471.530 2953.650 3474.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 -28.670 49.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 -28.670 229.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 -28.670 409.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 -28.670 589.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 -28.670 769.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 -28.670 949.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 -28.670 1129.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 -28.670 1669.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 -28.670 1849.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 -28.670 2029.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 -28.670 2209.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 -28.670 2389.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 -28.670 2569.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.170 -28.670 2749.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 236.240 49.270 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 236.240 229.270 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 236.240 409.270 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 236.240 589.270 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 236.240 1849.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 236.240 2029.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 236.240 2209.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 236.240 2389.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 236.240 2569.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.170 236.240 2749.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 1137.680 49.270 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 1137.680 229.270 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 1137.680 409.270 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 1137.680 589.270 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 236.240 769.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 236.240 949.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 236.240 1129.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 -28.670 1309.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 -28.670 1489.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 236.240 1669.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 1946.080 1849.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 1946.080 2029.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 1946.080 2209.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 2203.920 49.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 2203.920 229.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 2203.920 409.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 2203.920 589.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 3488.880 769.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 3488.880 949.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 3488.880 1129.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 3488.880 1309.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 3488.880 1489.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 3488.880 1669.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 3488.880 1849.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 3488.880 2029.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 3488.880 2209.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 1946.080 2389.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 1946.080 2569.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.170 1946.080 2749.270 3548.350 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 70.130 2963.250 73.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 250.130 2963.250 253.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 430.130 2963.250 433.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 610.130 2963.250 613.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 790.130 2963.250 793.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 970.130 2963.250 973.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1150.130 2963.250 1153.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1510.130 2963.250 1513.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1690.130 2963.250 1693.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2050.130 2963.250 2053.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2230.130 2963.250 2233.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2410.130 2963.250 2413.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2950.130 2963.250 2953.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3130.130 2963.250 3133.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 -38.270 67.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 -38.270 247.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 -38.270 427.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 -38.270 607.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 -38.270 787.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 -38.270 967.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 -38.270 1147.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 -38.270 1687.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 -38.270 1867.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 -38.270 2047.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 -38.270 2227.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 -38.270 2407.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 -38.270 2587.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2764.770 -38.270 2767.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 236.240 67.870 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 236.240 247.870 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 236.240 427.870 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 236.240 607.870 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 236.240 1867.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 236.240 2047.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 236.240 2227.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 236.240 2407.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 236.240 2587.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2764.770 236.240 2767.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 1137.680 67.870 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 1137.680 247.870 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 1137.680 427.870 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 1137.680 607.870 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 236.240 787.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 236.240 967.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 236.240 1147.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 -38.270 1327.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 -38.270 1507.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 236.240 1687.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 1946.080 1867.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 1946.080 2047.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 1946.080 2227.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 2203.920 67.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 2203.920 247.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 2203.920 427.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 2203.920 607.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 3488.880 787.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 3488.880 967.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 3488.880 1147.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 3488.880 1327.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 3488.880 1507.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 3488.880 1687.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 3488.880 1867.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 3488.880 2047.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 3488.880 2227.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 1946.080 2407.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 1946.080 2587.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2764.770 1946.080 2767.870 3557.950 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 141.530 2953.650 144.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 321.530 2953.650 324.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 501.530 2953.650 504.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 681.530 2953.650 684.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 861.530 2953.650 864.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1041.530 2953.650 1044.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1221.530 2953.650 1224.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1401.530 2953.650 1404.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1581.530 2953.650 1584.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1761.530 2953.650 1764.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1941.530 2953.650 1944.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2121.530 2953.650 2124.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2301.530 2953.650 2304.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2481.530 2953.650 2484.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2661.530 2953.650 2664.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2841.530 2953.650 2844.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3021.530 2953.650 3024.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3201.530 2953.650 3204.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3381.530 2953.650 3384.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.170 -28.670 139.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 -28.670 319.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 -28.670 499.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 -28.670 679.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 -28.670 859.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1036.170 -28.670 1039.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 -28.670 1219.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 -28.670 1759.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 -28.670 1939.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 -28.670 2119.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 -28.670 2299.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 -28.670 2479.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2656.170 -28.670 2659.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.170 -28.670 2839.270 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.170 236.240 139.270 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 236.240 319.270 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 236.240 499.270 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 236.240 679.270 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 236.240 1759.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 236.240 1939.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 236.240 2119.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 236.240 2299.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 236.240 2479.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2656.170 236.240 2659.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.170 236.240 2839.270 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.170 1137.680 139.270 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 1137.680 319.270 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 1137.680 499.270 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 1137.680 679.270 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 2203.920 679.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 236.240 859.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1036.170 236.240 1039.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 236.240 1219.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 -28.670 1399.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1576.170 -28.670 1579.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 1946.080 1759.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 1946.080 1939.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 1946.080 2119.270 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.170 2203.920 139.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 2203.920 319.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 2203.920 499.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 3488.880 679.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 3488.880 859.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1036.170 3488.880 1039.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 3488.880 1219.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 3488.880 1399.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1576.170 3488.880 1579.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 3488.880 1759.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 3488.880 1939.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 3488.880 2119.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 1946.080 2299.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 1946.080 2479.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2656.170 1946.080 2659.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.170 1946.080 2839.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 160.130 2963.250 163.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 340.130 2963.250 343.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 520.130 2963.250 523.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 700.130 2963.250 703.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 880.130 2963.250 883.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1060.130 2963.250 1063.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1240.130 2963.250 1243.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1420.130 2963.250 1423.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1600.130 2963.250 1603.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1780.130 2963.250 1783.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1960.130 2963.250 1963.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2140.130 2963.250 2143.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2320.130 2963.250 2323.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2500.130 2963.250 2503.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2680.130 2963.250 2683.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2860.130 2963.250 2863.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3040.130 2963.250 3043.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3220.130 2963.250 3223.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3400.130 2963.250 3403.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.770 -38.270 157.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 -38.270 337.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 -38.270 517.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 -38.270 697.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 -38.270 877.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.770 -38.270 1057.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 -38.270 1237.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 -38.270 1777.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 -38.270 1957.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 -38.270 2137.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 -38.270 2317.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 -38.270 2497.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2674.770 -38.270 2677.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.770 -38.270 2857.870 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.770 236.240 157.870 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 236.240 337.870 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 236.240 517.870 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 236.240 1777.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 236.240 1957.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 236.240 2137.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 236.240 2317.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 236.240 2497.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2674.770 236.240 2677.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.770 236.240 2857.870 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.770 1137.680 157.870 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 1137.680 337.870 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 1137.680 517.870 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 236.240 697.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 236.240 877.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.770 236.240 1057.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 236.240 1237.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 -38.270 1417.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 -38.270 1597.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 1946.080 1777.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 1946.080 1957.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 1946.080 2137.870 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.770 2203.920 157.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 2203.920 337.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 2203.920 517.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 3488.880 697.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 3488.880 877.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.770 3488.880 1057.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 3488.880 1237.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 3488.880 1417.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 3488.880 1597.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 3488.880 1777.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 3488.880 1957.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 3488.880 2137.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 1946.080 2317.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 1946.080 2497.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2674.770 1946.080 2677.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.770 1946.080 2857.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 104.090 2934.450 107.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 284.090 2934.450 287.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 464.090 2934.450 467.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 644.090 2934.450 647.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 824.090 2934.450 827.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1004.090 2934.450 1007.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1184.090 2934.450 1187.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1364.090 2934.450 1367.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1544.090 2934.450 1547.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1724.090 2934.450 1727.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1904.090 2934.450 1907.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2084.090 2934.450 2087.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2264.090 2934.450 2267.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2444.090 2934.450 2447.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2624.090 2934.450 2627.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2804.090 2934.450 2807.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2984.090 2934.450 2987.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3164.090 2934.450 3167.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3344.090 2934.450 3347.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 -9.470 102.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 -9.470 282.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 -9.470 462.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 -9.470 642.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 -9.470 822.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 -9.470 1002.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 -9.470 1182.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 -9.470 1722.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 -9.470 1902.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 -9.470 2082.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 -9.470 2262.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 -9.470 2442.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 -9.470 2622.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 -9.470 2802.070 31.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 236.000 102.070 517.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 236.000 282.070 517.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 236.000 462.070 517.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 236.000 642.070 517.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 236.000 1722.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 236.000 1902.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 236.000 2082.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 236.000 2262.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 236.000 2442.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 236.000 2622.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 236.000 2802.070 776.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 1137.440 102.070 1584.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 1137.440 282.070 1584.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1137.440 462.070 1584.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1137.440 642.070 1584.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2203.680 642.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 236.000 822.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 236.000 1002.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 236.000 1182.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 -9.470 1362.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 -9.470 1542.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 1945.840 1722.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 1945.840 1902.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 1945.840 2082.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 1945.840 2262.070 2481.760 ;
    END
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 2203.680 102.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 2203.680 282.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2203.680 462.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 3488.640 642.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 3488.640 822.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 3488.640 1002.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 3488.640 1182.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 3488.640 1362.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 3488.640 1542.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 3488.640 1722.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 3488.640 1902.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 3488.640 2082.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 3488.640 2262.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 1945.840 2442.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 1945.840 2622.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 1945.840 2802.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 122.930 2944.050 126.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 302.930 2944.050 306.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 482.930 2944.050 486.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 662.930 2944.050 666.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 842.930 2944.050 846.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1022.930 2944.050 1026.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1202.930 2944.050 1206.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1382.930 2944.050 1386.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1562.930 2944.050 1566.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1742.930 2944.050 1746.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1922.930 2944.050 1926.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2102.930 2944.050 2106.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2282.930 2944.050 2286.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2462.930 2944.050 2466.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2642.930 2944.050 2646.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2822.930 2944.050 2826.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3002.930 2944.050 3006.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3182.930 2944.050 3186.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3362.930 2944.050 3366.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.570 -19.070 120.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 -19.070 300.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 -19.070 480.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 -19.070 660.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 -19.070 840.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.570 -19.070 1020.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 -19.070 1200.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 -19.070 1740.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 -19.070 1920.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 -19.070 2100.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 -19.070 2280.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 -19.070 2460.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2637.570 -19.070 2640.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2817.570 -19.070 2820.670 30.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.570 236.240 120.670 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 236.240 300.670 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 236.240 480.670 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 236.240 660.670 517.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 236.240 1740.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 236.240 1920.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 236.240 2100.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 236.240 2280.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 236.240 2460.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2637.570 236.240 2640.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2817.570 236.240 2820.670 776.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.570 1137.680 120.670 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 1137.680 300.670 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 1137.680 480.670 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 1137.680 660.670 1583.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 2203.920 660.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 236.240 840.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.570 236.240 1020.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 236.240 1200.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 -19.070 1380.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.570 -19.070 1560.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 1946.080 1740.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 1946.080 1920.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 1946.080 2100.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 1946.080 2280.670 2481.520 ;
    END
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.570 2203.920 120.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 2203.920 300.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 2203.920 480.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 3488.880 660.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 3488.880 840.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.570 3488.880 1020.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 3488.880 1200.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 3488.880 1380.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.570 3488.880 1560.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 3488.880 1740.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 3488.880 1920.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 3488.880 2100.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 3488.880 2280.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 1946.080 2460.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2637.570 1946.080 2640.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2817.570 1946.080 2820.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2914.100 3508.885 ;
      LAYER met1 ;
        RECT 2.370 10.240 2917.250 3509.040 ;
      LAYER met2 ;
        RECT 2.390 3517.320 40.150 3518.050 ;
        RECT 41.270 3517.320 121.110 3518.050 ;
        RECT 122.230 3517.320 202.070 3518.050 ;
        RECT 203.190 3517.320 283.490 3518.050 ;
        RECT 284.610 3517.320 364.450 3518.050 ;
        RECT 365.570 3517.320 445.410 3518.050 ;
        RECT 446.530 3517.320 526.830 3518.050 ;
        RECT 527.950 3517.320 607.790 3518.050 ;
        RECT 608.910 3517.320 688.750 3518.050 ;
        RECT 689.870 3517.320 770.170 3518.050 ;
        RECT 771.290 3517.320 851.130 3518.050 ;
        RECT 852.250 3517.320 932.090 3518.050 ;
        RECT 933.210 3517.320 1013.510 3518.050 ;
        RECT 1014.630 3517.320 1094.470 3518.050 ;
        RECT 1095.590 3517.320 1175.430 3518.050 ;
        RECT 1176.550 3517.320 1256.850 3518.050 ;
        RECT 1257.970 3517.320 1337.810 3518.050 ;
        RECT 1338.930 3517.320 1418.770 3518.050 ;
        RECT 1419.890 3517.320 1500.190 3518.050 ;
        RECT 1501.310 3517.320 1581.150 3518.050 ;
        RECT 1582.270 3517.320 1662.110 3518.050 ;
        RECT 1663.230 3517.320 1743.530 3518.050 ;
        RECT 1744.650 3517.320 1824.490 3518.050 ;
        RECT 1825.610 3517.320 1905.450 3518.050 ;
        RECT 1906.570 3517.320 1986.870 3518.050 ;
        RECT 1987.990 3517.320 2067.830 3518.050 ;
        RECT 2068.950 3517.320 2148.790 3518.050 ;
        RECT 2149.910 3517.320 2230.210 3518.050 ;
        RECT 2231.330 3517.320 2311.170 3518.050 ;
        RECT 2312.290 3517.320 2392.130 3518.050 ;
        RECT 2393.250 3517.320 2473.550 3518.050 ;
        RECT 2474.670 3517.320 2554.510 3518.050 ;
        RECT 2555.630 3517.320 2635.470 3518.050 ;
        RECT 2636.590 3517.320 2716.890 3518.050 ;
        RECT 2718.010 3517.320 2797.850 3518.050 ;
        RECT 2798.970 3517.320 2878.810 3518.050 ;
        RECT 2879.930 3517.320 2917.220 3518.050 ;
        RECT 2.390 2.680 2917.220 3517.320 ;
        RECT 2.390 1.630 2.430 2.680 ;
        RECT 3.550 1.630 7.950 2.680 ;
        RECT 9.070 1.630 13.930 2.680 ;
        RECT 15.050 1.630 19.910 2.680 ;
        RECT 21.030 1.630 25.890 2.680 ;
        RECT 27.010 1.630 31.870 2.680 ;
        RECT 32.990 1.630 37.850 2.680 ;
        RECT 38.970 1.630 43.370 2.680 ;
        RECT 44.490 1.630 49.350 2.680 ;
        RECT 50.470 1.630 55.330 2.680 ;
        RECT 56.450 1.630 61.310 2.680 ;
        RECT 62.430 1.630 67.290 2.680 ;
        RECT 68.410 1.630 73.270 2.680 ;
        RECT 74.390 1.630 79.250 2.680 ;
        RECT 80.370 1.630 84.770 2.680 ;
        RECT 85.890 1.630 90.750 2.680 ;
        RECT 91.870 1.630 96.730 2.680 ;
        RECT 97.850 1.630 102.710 2.680 ;
        RECT 103.830 1.630 108.690 2.680 ;
        RECT 109.810 1.630 114.670 2.680 ;
        RECT 115.790 1.630 120.650 2.680 ;
        RECT 121.770 1.630 126.170 2.680 ;
        RECT 127.290 1.630 132.150 2.680 ;
        RECT 133.270 1.630 138.130 2.680 ;
        RECT 139.250 1.630 144.110 2.680 ;
        RECT 145.230 1.630 150.090 2.680 ;
        RECT 151.210 1.630 156.070 2.680 ;
        RECT 157.190 1.630 161.590 2.680 ;
        RECT 162.710 1.630 167.570 2.680 ;
        RECT 168.690 1.630 173.550 2.680 ;
        RECT 174.670 1.630 179.530 2.680 ;
        RECT 180.650 1.630 185.510 2.680 ;
        RECT 186.630 1.630 191.490 2.680 ;
        RECT 192.610 1.630 197.470 2.680 ;
        RECT 198.590 1.630 202.990 2.680 ;
        RECT 204.110 1.630 208.970 2.680 ;
        RECT 210.090 1.630 214.950 2.680 ;
        RECT 216.070 1.630 220.930 2.680 ;
        RECT 222.050 1.630 226.910 2.680 ;
        RECT 228.030 1.630 232.890 2.680 ;
        RECT 234.010 1.630 238.870 2.680 ;
        RECT 239.990 1.630 244.390 2.680 ;
        RECT 245.510 1.630 250.370 2.680 ;
        RECT 251.490 1.630 256.350 2.680 ;
        RECT 257.470 1.630 262.330 2.680 ;
        RECT 263.450 1.630 268.310 2.680 ;
        RECT 269.430 1.630 274.290 2.680 ;
        RECT 275.410 1.630 279.810 2.680 ;
        RECT 280.930 1.630 285.790 2.680 ;
        RECT 286.910 1.630 291.770 2.680 ;
        RECT 292.890 1.630 297.750 2.680 ;
        RECT 298.870 1.630 303.730 2.680 ;
        RECT 304.850 1.630 309.710 2.680 ;
        RECT 310.830 1.630 315.690 2.680 ;
        RECT 316.810 1.630 321.210 2.680 ;
        RECT 322.330 1.630 327.190 2.680 ;
        RECT 328.310 1.630 333.170 2.680 ;
        RECT 334.290 1.630 339.150 2.680 ;
        RECT 340.270 1.630 345.130 2.680 ;
        RECT 346.250 1.630 351.110 2.680 ;
        RECT 352.230 1.630 357.090 2.680 ;
        RECT 358.210 1.630 362.610 2.680 ;
        RECT 363.730 1.630 368.590 2.680 ;
        RECT 369.710 1.630 374.570 2.680 ;
        RECT 375.690 1.630 380.550 2.680 ;
        RECT 381.670 1.630 386.530 2.680 ;
        RECT 387.650 1.630 392.510 2.680 ;
        RECT 393.630 1.630 398.030 2.680 ;
        RECT 399.150 1.630 404.010 2.680 ;
        RECT 405.130 1.630 409.990 2.680 ;
        RECT 411.110 1.630 415.970 2.680 ;
        RECT 417.090 1.630 421.950 2.680 ;
        RECT 423.070 1.630 427.930 2.680 ;
        RECT 429.050 1.630 433.910 2.680 ;
        RECT 435.030 1.630 439.430 2.680 ;
        RECT 440.550 1.630 445.410 2.680 ;
        RECT 446.530 1.630 451.390 2.680 ;
        RECT 452.510 1.630 457.370 2.680 ;
        RECT 458.490 1.630 463.350 2.680 ;
        RECT 464.470 1.630 469.330 2.680 ;
        RECT 470.450 1.630 475.310 2.680 ;
        RECT 476.430 1.630 480.830 2.680 ;
        RECT 481.950 1.630 486.810 2.680 ;
        RECT 487.930 1.630 492.790 2.680 ;
        RECT 493.910 1.630 498.770 2.680 ;
        RECT 499.890 1.630 504.750 2.680 ;
        RECT 505.870 1.630 510.730 2.680 ;
        RECT 511.850 1.630 516.250 2.680 ;
        RECT 517.370 1.630 522.230 2.680 ;
        RECT 523.350 1.630 528.210 2.680 ;
        RECT 529.330 1.630 534.190 2.680 ;
        RECT 535.310 1.630 540.170 2.680 ;
        RECT 541.290 1.630 546.150 2.680 ;
        RECT 547.270 1.630 552.130 2.680 ;
        RECT 553.250 1.630 557.650 2.680 ;
        RECT 558.770 1.630 563.630 2.680 ;
        RECT 564.750 1.630 569.610 2.680 ;
        RECT 570.730 1.630 575.590 2.680 ;
        RECT 576.710 1.630 581.570 2.680 ;
        RECT 582.690 1.630 587.550 2.680 ;
        RECT 588.670 1.630 593.530 2.680 ;
        RECT 594.650 1.630 599.050 2.680 ;
        RECT 600.170 1.630 605.030 2.680 ;
        RECT 606.150 1.630 611.010 2.680 ;
        RECT 612.130 1.630 616.990 2.680 ;
        RECT 618.110 1.630 622.970 2.680 ;
        RECT 624.090 1.630 628.950 2.680 ;
        RECT 630.070 1.630 634.470 2.680 ;
        RECT 635.590 1.630 640.450 2.680 ;
        RECT 641.570 1.630 646.430 2.680 ;
        RECT 647.550 1.630 652.410 2.680 ;
        RECT 653.530 1.630 658.390 2.680 ;
        RECT 659.510 1.630 664.370 2.680 ;
        RECT 665.490 1.630 670.350 2.680 ;
        RECT 671.470 1.630 675.870 2.680 ;
        RECT 676.990 1.630 681.850 2.680 ;
        RECT 682.970 1.630 687.830 2.680 ;
        RECT 688.950 1.630 693.810 2.680 ;
        RECT 694.930 1.630 699.790 2.680 ;
        RECT 700.910 1.630 705.770 2.680 ;
        RECT 706.890 1.630 711.750 2.680 ;
        RECT 712.870 1.630 717.270 2.680 ;
        RECT 718.390 1.630 723.250 2.680 ;
        RECT 724.370 1.630 729.230 2.680 ;
        RECT 730.350 1.630 735.210 2.680 ;
        RECT 736.330 1.630 741.190 2.680 ;
        RECT 742.310 1.630 747.170 2.680 ;
        RECT 748.290 1.630 752.690 2.680 ;
        RECT 753.810 1.630 758.670 2.680 ;
        RECT 759.790 1.630 764.650 2.680 ;
        RECT 765.770 1.630 770.630 2.680 ;
        RECT 771.750 1.630 776.610 2.680 ;
        RECT 777.730 1.630 782.590 2.680 ;
        RECT 783.710 1.630 788.570 2.680 ;
        RECT 789.690 1.630 794.090 2.680 ;
        RECT 795.210 1.630 800.070 2.680 ;
        RECT 801.190 1.630 806.050 2.680 ;
        RECT 807.170 1.630 812.030 2.680 ;
        RECT 813.150 1.630 818.010 2.680 ;
        RECT 819.130 1.630 823.990 2.680 ;
        RECT 825.110 1.630 829.970 2.680 ;
        RECT 831.090 1.630 835.490 2.680 ;
        RECT 836.610 1.630 841.470 2.680 ;
        RECT 842.590 1.630 847.450 2.680 ;
        RECT 848.570 1.630 853.430 2.680 ;
        RECT 854.550 1.630 859.410 2.680 ;
        RECT 860.530 1.630 865.390 2.680 ;
        RECT 866.510 1.630 870.910 2.680 ;
        RECT 872.030 1.630 876.890 2.680 ;
        RECT 878.010 1.630 882.870 2.680 ;
        RECT 883.990 1.630 888.850 2.680 ;
        RECT 889.970 1.630 894.830 2.680 ;
        RECT 895.950 1.630 900.810 2.680 ;
        RECT 901.930 1.630 906.790 2.680 ;
        RECT 907.910 1.630 912.310 2.680 ;
        RECT 913.430 1.630 918.290 2.680 ;
        RECT 919.410 1.630 924.270 2.680 ;
        RECT 925.390 1.630 930.250 2.680 ;
        RECT 931.370 1.630 936.230 2.680 ;
        RECT 937.350 1.630 942.210 2.680 ;
        RECT 943.330 1.630 948.190 2.680 ;
        RECT 949.310 1.630 953.710 2.680 ;
        RECT 954.830 1.630 959.690 2.680 ;
        RECT 960.810 1.630 965.670 2.680 ;
        RECT 966.790 1.630 971.650 2.680 ;
        RECT 972.770 1.630 977.630 2.680 ;
        RECT 978.750 1.630 983.610 2.680 ;
        RECT 984.730 1.630 989.130 2.680 ;
        RECT 990.250 1.630 995.110 2.680 ;
        RECT 996.230 1.630 1001.090 2.680 ;
        RECT 1002.210 1.630 1007.070 2.680 ;
        RECT 1008.190 1.630 1013.050 2.680 ;
        RECT 1014.170 1.630 1019.030 2.680 ;
        RECT 1020.150 1.630 1025.010 2.680 ;
        RECT 1026.130 1.630 1030.530 2.680 ;
        RECT 1031.650 1.630 1036.510 2.680 ;
        RECT 1037.630 1.630 1042.490 2.680 ;
        RECT 1043.610 1.630 1048.470 2.680 ;
        RECT 1049.590 1.630 1054.450 2.680 ;
        RECT 1055.570 1.630 1060.430 2.680 ;
        RECT 1061.550 1.630 1066.410 2.680 ;
        RECT 1067.530 1.630 1071.930 2.680 ;
        RECT 1073.050 1.630 1077.910 2.680 ;
        RECT 1079.030 1.630 1083.890 2.680 ;
        RECT 1085.010 1.630 1089.870 2.680 ;
        RECT 1090.990 1.630 1095.850 2.680 ;
        RECT 1096.970 1.630 1101.830 2.680 ;
        RECT 1102.950 1.630 1107.350 2.680 ;
        RECT 1108.470 1.630 1113.330 2.680 ;
        RECT 1114.450 1.630 1119.310 2.680 ;
        RECT 1120.430 1.630 1125.290 2.680 ;
        RECT 1126.410 1.630 1131.270 2.680 ;
        RECT 1132.390 1.630 1137.250 2.680 ;
        RECT 1138.370 1.630 1143.230 2.680 ;
        RECT 1144.350 1.630 1148.750 2.680 ;
        RECT 1149.870 1.630 1154.730 2.680 ;
        RECT 1155.850 1.630 1160.710 2.680 ;
        RECT 1161.830 1.630 1166.690 2.680 ;
        RECT 1167.810 1.630 1172.670 2.680 ;
        RECT 1173.790 1.630 1178.650 2.680 ;
        RECT 1179.770 1.630 1184.630 2.680 ;
        RECT 1185.750 1.630 1190.150 2.680 ;
        RECT 1191.270 1.630 1196.130 2.680 ;
        RECT 1197.250 1.630 1202.110 2.680 ;
        RECT 1203.230 1.630 1208.090 2.680 ;
        RECT 1209.210 1.630 1214.070 2.680 ;
        RECT 1215.190 1.630 1220.050 2.680 ;
        RECT 1221.170 1.630 1225.570 2.680 ;
        RECT 1226.690 1.630 1231.550 2.680 ;
        RECT 1232.670 1.630 1237.530 2.680 ;
        RECT 1238.650 1.630 1243.510 2.680 ;
        RECT 1244.630 1.630 1249.490 2.680 ;
        RECT 1250.610 1.630 1255.470 2.680 ;
        RECT 1256.590 1.630 1261.450 2.680 ;
        RECT 1262.570 1.630 1266.970 2.680 ;
        RECT 1268.090 1.630 1272.950 2.680 ;
        RECT 1274.070 1.630 1278.930 2.680 ;
        RECT 1280.050 1.630 1284.910 2.680 ;
        RECT 1286.030 1.630 1290.890 2.680 ;
        RECT 1292.010 1.630 1296.870 2.680 ;
        RECT 1297.990 1.630 1302.850 2.680 ;
        RECT 1303.970 1.630 1308.370 2.680 ;
        RECT 1309.490 1.630 1314.350 2.680 ;
        RECT 1315.470 1.630 1320.330 2.680 ;
        RECT 1321.450 1.630 1326.310 2.680 ;
        RECT 1327.430 1.630 1332.290 2.680 ;
        RECT 1333.410 1.630 1338.270 2.680 ;
        RECT 1339.390 1.630 1343.790 2.680 ;
        RECT 1344.910 1.630 1349.770 2.680 ;
        RECT 1350.890 1.630 1355.750 2.680 ;
        RECT 1356.870 1.630 1361.730 2.680 ;
        RECT 1362.850 1.630 1367.710 2.680 ;
        RECT 1368.830 1.630 1373.690 2.680 ;
        RECT 1374.810 1.630 1379.670 2.680 ;
        RECT 1380.790 1.630 1385.190 2.680 ;
        RECT 1386.310 1.630 1391.170 2.680 ;
        RECT 1392.290 1.630 1397.150 2.680 ;
        RECT 1398.270 1.630 1403.130 2.680 ;
        RECT 1404.250 1.630 1409.110 2.680 ;
        RECT 1410.230 1.630 1415.090 2.680 ;
        RECT 1416.210 1.630 1421.070 2.680 ;
        RECT 1422.190 1.630 1426.590 2.680 ;
        RECT 1427.710 1.630 1432.570 2.680 ;
        RECT 1433.690 1.630 1438.550 2.680 ;
        RECT 1439.670 1.630 1444.530 2.680 ;
        RECT 1445.650 1.630 1450.510 2.680 ;
        RECT 1451.630 1.630 1456.490 2.680 ;
        RECT 1457.610 1.630 1462.470 2.680 ;
        RECT 1463.590 1.630 1467.990 2.680 ;
        RECT 1469.110 1.630 1473.970 2.680 ;
        RECT 1475.090 1.630 1479.950 2.680 ;
        RECT 1481.070 1.630 1485.930 2.680 ;
        RECT 1487.050 1.630 1491.910 2.680 ;
        RECT 1493.030 1.630 1497.890 2.680 ;
        RECT 1499.010 1.630 1503.410 2.680 ;
        RECT 1504.530 1.630 1509.390 2.680 ;
        RECT 1510.510 1.630 1515.370 2.680 ;
        RECT 1516.490 1.630 1521.350 2.680 ;
        RECT 1522.470 1.630 1527.330 2.680 ;
        RECT 1528.450 1.630 1533.310 2.680 ;
        RECT 1534.430 1.630 1539.290 2.680 ;
        RECT 1540.410 1.630 1544.810 2.680 ;
        RECT 1545.930 1.630 1550.790 2.680 ;
        RECT 1551.910 1.630 1556.770 2.680 ;
        RECT 1557.890 1.630 1562.750 2.680 ;
        RECT 1563.870 1.630 1568.730 2.680 ;
        RECT 1569.850 1.630 1574.710 2.680 ;
        RECT 1575.830 1.630 1580.690 2.680 ;
        RECT 1581.810 1.630 1586.210 2.680 ;
        RECT 1587.330 1.630 1592.190 2.680 ;
        RECT 1593.310 1.630 1598.170 2.680 ;
        RECT 1599.290 1.630 1604.150 2.680 ;
        RECT 1605.270 1.630 1610.130 2.680 ;
        RECT 1611.250 1.630 1616.110 2.680 ;
        RECT 1617.230 1.630 1621.630 2.680 ;
        RECT 1622.750 1.630 1627.610 2.680 ;
        RECT 1628.730 1.630 1633.590 2.680 ;
        RECT 1634.710 1.630 1639.570 2.680 ;
        RECT 1640.690 1.630 1645.550 2.680 ;
        RECT 1646.670 1.630 1651.530 2.680 ;
        RECT 1652.650 1.630 1657.510 2.680 ;
        RECT 1658.630 1.630 1663.030 2.680 ;
        RECT 1664.150 1.630 1669.010 2.680 ;
        RECT 1670.130 1.630 1674.990 2.680 ;
        RECT 1676.110 1.630 1680.970 2.680 ;
        RECT 1682.090 1.630 1686.950 2.680 ;
        RECT 1688.070 1.630 1692.930 2.680 ;
        RECT 1694.050 1.630 1698.910 2.680 ;
        RECT 1700.030 1.630 1704.430 2.680 ;
        RECT 1705.550 1.630 1710.410 2.680 ;
        RECT 1711.530 1.630 1716.390 2.680 ;
        RECT 1717.510 1.630 1722.370 2.680 ;
        RECT 1723.490 1.630 1728.350 2.680 ;
        RECT 1729.470 1.630 1734.330 2.680 ;
        RECT 1735.450 1.630 1739.850 2.680 ;
        RECT 1740.970 1.630 1745.830 2.680 ;
        RECT 1746.950 1.630 1751.810 2.680 ;
        RECT 1752.930 1.630 1757.790 2.680 ;
        RECT 1758.910 1.630 1763.770 2.680 ;
        RECT 1764.890 1.630 1769.750 2.680 ;
        RECT 1770.870 1.630 1775.730 2.680 ;
        RECT 1776.850 1.630 1781.250 2.680 ;
        RECT 1782.370 1.630 1787.230 2.680 ;
        RECT 1788.350 1.630 1793.210 2.680 ;
        RECT 1794.330 1.630 1799.190 2.680 ;
        RECT 1800.310 1.630 1805.170 2.680 ;
        RECT 1806.290 1.630 1811.150 2.680 ;
        RECT 1812.270 1.630 1817.130 2.680 ;
        RECT 1818.250 1.630 1822.650 2.680 ;
        RECT 1823.770 1.630 1828.630 2.680 ;
        RECT 1829.750 1.630 1834.610 2.680 ;
        RECT 1835.730 1.630 1840.590 2.680 ;
        RECT 1841.710 1.630 1846.570 2.680 ;
        RECT 1847.690 1.630 1852.550 2.680 ;
        RECT 1853.670 1.630 1858.070 2.680 ;
        RECT 1859.190 1.630 1864.050 2.680 ;
        RECT 1865.170 1.630 1870.030 2.680 ;
        RECT 1871.150 1.630 1876.010 2.680 ;
        RECT 1877.130 1.630 1881.990 2.680 ;
        RECT 1883.110 1.630 1887.970 2.680 ;
        RECT 1889.090 1.630 1893.950 2.680 ;
        RECT 1895.070 1.630 1899.470 2.680 ;
        RECT 1900.590 1.630 1905.450 2.680 ;
        RECT 1906.570 1.630 1911.430 2.680 ;
        RECT 1912.550 1.630 1917.410 2.680 ;
        RECT 1918.530 1.630 1923.390 2.680 ;
        RECT 1924.510 1.630 1929.370 2.680 ;
        RECT 1930.490 1.630 1935.350 2.680 ;
        RECT 1936.470 1.630 1940.870 2.680 ;
        RECT 1941.990 1.630 1946.850 2.680 ;
        RECT 1947.970 1.630 1952.830 2.680 ;
        RECT 1953.950 1.630 1958.810 2.680 ;
        RECT 1959.930 1.630 1964.790 2.680 ;
        RECT 1965.910 1.630 1970.770 2.680 ;
        RECT 1971.890 1.630 1976.290 2.680 ;
        RECT 1977.410 1.630 1982.270 2.680 ;
        RECT 1983.390 1.630 1988.250 2.680 ;
        RECT 1989.370 1.630 1994.230 2.680 ;
        RECT 1995.350 1.630 2000.210 2.680 ;
        RECT 2001.330 1.630 2006.190 2.680 ;
        RECT 2007.310 1.630 2012.170 2.680 ;
        RECT 2013.290 1.630 2017.690 2.680 ;
        RECT 2018.810 1.630 2023.670 2.680 ;
        RECT 2024.790 1.630 2029.650 2.680 ;
        RECT 2030.770 1.630 2035.630 2.680 ;
        RECT 2036.750 1.630 2041.610 2.680 ;
        RECT 2042.730 1.630 2047.590 2.680 ;
        RECT 2048.710 1.630 2053.570 2.680 ;
        RECT 2054.690 1.630 2059.090 2.680 ;
        RECT 2060.210 1.630 2065.070 2.680 ;
        RECT 2066.190 1.630 2071.050 2.680 ;
        RECT 2072.170 1.630 2077.030 2.680 ;
        RECT 2078.150 1.630 2083.010 2.680 ;
        RECT 2084.130 1.630 2088.990 2.680 ;
        RECT 2090.110 1.630 2094.510 2.680 ;
        RECT 2095.630 1.630 2100.490 2.680 ;
        RECT 2101.610 1.630 2106.470 2.680 ;
        RECT 2107.590 1.630 2112.450 2.680 ;
        RECT 2113.570 1.630 2118.430 2.680 ;
        RECT 2119.550 1.630 2124.410 2.680 ;
        RECT 2125.530 1.630 2130.390 2.680 ;
        RECT 2131.510 1.630 2135.910 2.680 ;
        RECT 2137.030 1.630 2141.890 2.680 ;
        RECT 2143.010 1.630 2147.870 2.680 ;
        RECT 2148.990 1.630 2153.850 2.680 ;
        RECT 2154.970 1.630 2159.830 2.680 ;
        RECT 2160.950 1.630 2165.810 2.680 ;
        RECT 2166.930 1.630 2171.790 2.680 ;
        RECT 2172.910 1.630 2177.310 2.680 ;
        RECT 2178.430 1.630 2183.290 2.680 ;
        RECT 2184.410 1.630 2189.270 2.680 ;
        RECT 2190.390 1.630 2195.250 2.680 ;
        RECT 2196.370 1.630 2201.230 2.680 ;
        RECT 2202.350 1.630 2207.210 2.680 ;
        RECT 2208.330 1.630 2212.730 2.680 ;
        RECT 2213.850 1.630 2218.710 2.680 ;
        RECT 2219.830 1.630 2224.690 2.680 ;
        RECT 2225.810 1.630 2230.670 2.680 ;
        RECT 2231.790 1.630 2236.650 2.680 ;
        RECT 2237.770 1.630 2242.630 2.680 ;
        RECT 2243.750 1.630 2248.610 2.680 ;
        RECT 2249.730 1.630 2254.130 2.680 ;
        RECT 2255.250 1.630 2260.110 2.680 ;
        RECT 2261.230 1.630 2266.090 2.680 ;
        RECT 2267.210 1.630 2272.070 2.680 ;
        RECT 2273.190 1.630 2278.050 2.680 ;
        RECT 2279.170 1.630 2284.030 2.680 ;
        RECT 2285.150 1.630 2290.010 2.680 ;
        RECT 2291.130 1.630 2295.530 2.680 ;
        RECT 2296.650 1.630 2301.510 2.680 ;
        RECT 2302.630 1.630 2307.490 2.680 ;
        RECT 2308.610 1.630 2313.470 2.680 ;
        RECT 2314.590 1.630 2319.450 2.680 ;
        RECT 2320.570 1.630 2325.430 2.680 ;
        RECT 2326.550 1.630 2330.950 2.680 ;
        RECT 2332.070 1.630 2336.930 2.680 ;
        RECT 2338.050 1.630 2342.910 2.680 ;
        RECT 2344.030 1.630 2348.890 2.680 ;
        RECT 2350.010 1.630 2354.870 2.680 ;
        RECT 2355.990 1.630 2360.850 2.680 ;
        RECT 2361.970 1.630 2366.830 2.680 ;
        RECT 2367.950 1.630 2372.350 2.680 ;
        RECT 2373.470 1.630 2378.330 2.680 ;
        RECT 2379.450 1.630 2384.310 2.680 ;
        RECT 2385.430 1.630 2390.290 2.680 ;
        RECT 2391.410 1.630 2396.270 2.680 ;
        RECT 2397.390 1.630 2402.250 2.680 ;
        RECT 2403.370 1.630 2408.230 2.680 ;
        RECT 2409.350 1.630 2413.750 2.680 ;
        RECT 2414.870 1.630 2419.730 2.680 ;
        RECT 2420.850 1.630 2425.710 2.680 ;
        RECT 2426.830 1.630 2431.690 2.680 ;
        RECT 2432.810 1.630 2437.670 2.680 ;
        RECT 2438.790 1.630 2443.650 2.680 ;
        RECT 2444.770 1.630 2449.170 2.680 ;
        RECT 2450.290 1.630 2455.150 2.680 ;
        RECT 2456.270 1.630 2461.130 2.680 ;
        RECT 2462.250 1.630 2467.110 2.680 ;
        RECT 2468.230 1.630 2473.090 2.680 ;
        RECT 2474.210 1.630 2479.070 2.680 ;
        RECT 2480.190 1.630 2485.050 2.680 ;
        RECT 2486.170 1.630 2490.570 2.680 ;
        RECT 2491.690 1.630 2496.550 2.680 ;
        RECT 2497.670 1.630 2502.530 2.680 ;
        RECT 2503.650 1.630 2508.510 2.680 ;
        RECT 2509.630 1.630 2514.490 2.680 ;
        RECT 2515.610 1.630 2520.470 2.680 ;
        RECT 2521.590 1.630 2526.450 2.680 ;
        RECT 2527.570 1.630 2531.970 2.680 ;
        RECT 2533.090 1.630 2537.950 2.680 ;
        RECT 2539.070 1.630 2543.930 2.680 ;
        RECT 2545.050 1.630 2549.910 2.680 ;
        RECT 2551.030 1.630 2555.890 2.680 ;
        RECT 2557.010 1.630 2561.870 2.680 ;
        RECT 2562.990 1.630 2567.390 2.680 ;
        RECT 2568.510 1.630 2573.370 2.680 ;
        RECT 2574.490 1.630 2579.350 2.680 ;
        RECT 2580.470 1.630 2585.330 2.680 ;
        RECT 2586.450 1.630 2591.310 2.680 ;
        RECT 2592.430 1.630 2597.290 2.680 ;
        RECT 2598.410 1.630 2603.270 2.680 ;
        RECT 2604.390 1.630 2608.790 2.680 ;
        RECT 2609.910 1.630 2614.770 2.680 ;
        RECT 2615.890 1.630 2620.750 2.680 ;
        RECT 2621.870 1.630 2626.730 2.680 ;
        RECT 2627.850 1.630 2632.710 2.680 ;
        RECT 2633.830 1.630 2638.690 2.680 ;
        RECT 2639.810 1.630 2644.670 2.680 ;
        RECT 2645.790 1.630 2650.190 2.680 ;
        RECT 2651.310 1.630 2656.170 2.680 ;
        RECT 2657.290 1.630 2662.150 2.680 ;
        RECT 2663.270 1.630 2668.130 2.680 ;
        RECT 2669.250 1.630 2674.110 2.680 ;
        RECT 2675.230 1.630 2680.090 2.680 ;
        RECT 2681.210 1.630 2685.610 2.680 ;
        RECT 2686.730 1.630 2691.590 2.680 ;
        RECT 2692.710 1.630 2697.570 2.680 ;
        RECT 2698.690 1.630 2703.550 2.680 ;
        RECT 2704.670 1.630 2709.530 2.680 ;
        RECT 2710.650 1.630 2715.510 2.680 ;
        RECT 2716.630 1.630 2721.490 2.680 ;
        RECT 2722.610 1.630 2727.010 2.680 ;
        RECT 2728.130 1.630 2732.990 2.680 ;
        RECT 2734.110 1.630 2738.970 2.680 ;
        RECT 2740.090 1.630 2744.950 2.680 ;
        RECT 2746.070 1.630 2750.930 2.680 ;
        RECT 2752.050 1.630 2756.910 2.680 ;
        RECT 2758.030 1.630 2762.890 2.680 ;
        RECT 2764.010 1.630 2768.410 2.680 ;
        RECT 2769.530 1.630 2774.390 2.680 ;
        RECT 2775.510 1.630 2780.370 2.680 ;
        RECT 2781.490 1.630 2786.350 2.680 ;
        RECT 2787.470 1.630 2792.330 2.680 ;
        RECT 2793.450 1.630 2798.310 2.680 ;
        RECT 2799.430 1.630 2803.830 2.680 ;
        RECT 2804.950 1.630 2809.810 2.680 ;
        RECT 2810.930 1.630 2815.790 2.680 ;
        RECT 2816.910 1.630 2821.770 2.680 ;
        RECT 2822.890 1.630 2827.750 2.680 ;
        RECT 2828.870 1.630 2833.730 2.680 ;
        RECT 2834.850 1.630 2839.710 2.680 ;
        RECT 2840.830 1.630 2845.230 2.680 ;
        RECT 2846.350 1.630 2851.210 2.680 ;
        RECT 2852.330 1.630 2857.190 2.680 ;
        RECT 2858.310 1.630 2863.170 2.680 ;
        RECT 2864.290 1.630 2869.150 2.680 ;
        RECT 2870.270 1.630 2875.130 2.680 ;
        RECT 2876.250 1.630 2881.110 2.680 ;
        RECT 2882.230 1.630 2886.630 2.680 ;
        RECT 2887.750 1.630 2892.610 2.680 ;
        RECT 2893.730 1.630 2898.590 2.680 ;
        RECT 2899.710 1.630 2904.570 2.680 ;
        RECT 2905.690 1.630 2910.550 2.680 ;
        RECT 2911.670 1.630 2916.530 2.680 ;
      LAYER met3 ;
        RECT 2.365 3487.700 2917.600 3508.965 ;
        RECT 2.800 3487.020 2917.600 3487.700 ;
        RECT 2.800 3485.700 2917.200 3487.020 ;
        RECT 2.365 3485.020 2917.200 3485.700 ;
        RECT 2.365 3422.420 2917.600 3485.020 ;
        RECT 2.800 3420.420 2917.600 3422.420 ;
        RECT 2.365 3420.380 2917.600 3420.420 ;
        RECT 2.365 3418.380 2917.200 3420.380 ;
        RECT 2.365 3357.140 2917.600 3418.380 ;
        RECT 2.800 3355.140 2917.600 3357.140 ;
        RECT 2.365 3354.420 2917.600 3355.140 ;
        RECT 2.365 3352.420 2917.200 3354.420 ;
        RECT 2.365 3291.860 2917.600 3352.420 ;
        RECT 2.800 3289.860 2917.600 3291.860 ;
        RECT 2.365 3287.780 2917.600 3289.860 ;
        RECT 2.365 3285.780 2917.200 3287.780 ;
        RECT 2.365 3226.580 2917.600 3285.780 ;
        RECT 2.800 3224.580 2917.600 3226.580 ;
        RECT 2.365 3221.140 2917.600 3224.580 ;
        RECT 2.365 3219.140 2917.200 3221.140 ;
        RECT 2.365 3161.300 2917.600 3219.140 ;
        RECT 2.800 3159.300 2917.600 3161.300 ;
        RECT 2.365 3155.180 2917.600 3159.300 ;
        RECT 2.365 3153.180 2917.200 3155.180 ;
        RECT 2.365 3096.700 2917.600 3153.180 ;
        RECT 2.800 3094.700 2917.600 3096.700 ;
        RECT 2.365 3088.540 2917.600 3094.700 ;
        RECT 2.365 3086.540 2917.200 3088.540 ;
        RECT 2.365 3031.420 2917.600 3086.540 ;
        RECT 2.800 3029.420 2917.600 3031.420 ;
        RECT 2.365 3021.900 2917.600 3029.420 ;
        RECT 2.365 3019.900 2917.200 3021.900 ;
        RECT 2.365 2966.140 2917.600 3019.900 ;
        RECT 2.800 2964.140 2917.600 2966.140 ;
        RECT 2.365 2955.940 2917.600 2964.140 ;
        RECT 2.365 2953.940 2917.200 2955.940 ;
        RECT 2.365 2900.860 2917.600 2953.940 ;
        RECT 2.800 2898.860 2917.600 2900.860 ;
        RECT 2.365 2889.300 2917.600 2898.860 ;
        RECT 2.365 2887.300 2917.200 2889.300 ;
        RECT 2.365 2835.580 2917.600 2887.300 ;
        RECT 2.800 2833.580 2917.600 2835.580 ;
        RECT 2.365 2822.660 2917.600 2833.580 ;
        RECT 2.365 2820.660 2917.200 2822.660 ;
        RECT 2.365 2770.300 2917.600 2820.660 ;
        RECT 2.800 2768.300 2917.600 2770.300 ;
        RECT 2.365 2756.700 2917.600 2768.300 ;
        RECT 2.365 2754.700 2917.200 2756.700 ;
        RECT 2.365 2705.020 2917.600 2754.700 ;
        RECT 2.800 2703.020 2917.600 2705.020 ;
        RECT 2.365 2690.060 2917.600 2703.020 ;
        RECT 2.365 2688.060 2917.200 2690.060 ;
        RECT 2.365 2640.420 2917.600 2688.060 ;
        RECT 2.800 2638.420 2917.600 2640.420 ;
        RECT 2.365 2623.420 2917.600 2638.420 ;
        RECT 2.365 2621.420 2917.200 2623.420 ;
        RECT 2.365 2575.140 2917.600 2621.420 ;
        RECT 2.800 2573.140 2917.600 2575.140 ;
        RECT 2.365 2557.460 2917.600 2573.140 ;
        RECT 2.365 2555.460 2917.200 2557.460 ;
        RECT 2.365 2509.860 2917.600 2555.460 ;
        RECT 2.800 2507.860 2917.600 2509.860 ;
        RECT 2.365 2490.820 2917.600 2507.860 ;
        RECT 2.365 2488.820 2917.200 2490.820 ;
        RECT 2.365 2444.580 2917.600 2488.820 ;
        RECT 2.800 2442.580 2917.600 2444.580 ;
        RECT 2.365 2424.180 2917.600 2442.580 ;
        RECT 2.365 2422.180 2917.200 2424.180 ;
        RECT 2.365 2379.300 2917.600 2422.180 ;
        RECT 2.800 2377.300 2917.600 2379.300 ;
        RECT 2.365 2358.220 2917.600 2377.300 ;
        RECT 2.365 2356.220 2917.200 2358.220 ;
        RECT 2.365 2314.020 2917.600 2356.220 ;
        RECT 2.800 2312.020 2917.600 2314.020 ;
        RECT 2.365 2291.580 2917.600 2312.020 ;
        RECT 2.365 2289.580 2917.200 2291.580 ;
        RECT 2.365 2248.740 2917.600 2289.580 ;
        RECT 2.800 2246.740 2917.600 2248.740 ;
        RECT 2.365 2224.940 2917.600 2246.740 ;
        RECT 2.365 2222.940 2917.200 2224.940 ;
        RECT 2.365 2184.140 2917.600 2222.940 ;
        RECT 2.800 2182.140 2917.600 2184.140 ;
        RECT 2.365 2158.980 2917.600 2182.140 ;
        RECT 2.365 2156.980 2917.200 2158.980 ;
        RECT 2.365 2118.860 2917.600 2156.980 ;
        RECT 2.800 2116.860 2917.600 2118.860 ;
        RECT 2.365 2092.340 2917.600 2116.860 ;
        RECT 2.365 2090.340 2917.200 2092.340 ;
        RECT 2.365 2053.580 2917.600 2090.340 ;
        RECT 2.800 2051.580 2917.600 2053.580 ;
        RECT 2.365 2025.700 2917.600 2051.580 ;
        RECT 2.365 2023.700 2917.200 2025.700 ;
        RECT 2.365 1988.300 2917.600 2023.700 ;
        RECT 2.800 1986.300 2917.600 1988.300 ;
        RECT 2.365 1959.740 2917.600 1986.300 ;
        RECT 2.365 1957.740 2917.200 1959.740 ;
        RECT 2.365 1923.020 2917.600 1957.740 ;
        RECT 2.800 1921.020 2917.600 1923.020 ;
        RECT 2.365 1893.100 2917.600 1921.020 ;
        RECT 2.365 1891.100 2917.200 1893.100 ;
        RECT 2.365 1857.740 2917.600 1891.100 ;
        RECT 2.800 1855.740 2917.600 1857.740 ;
        RECT 2.365 1826.460 2917.600 1855.740 ;
        RECT 2.365 1824.460 2917.200 1826.460 ;
        RECT 2.365 1793.140 2917.600 1824.460 ;
        RECT 2.800 1791.140 2917.600 1793.140 ;
        RECT 2.365 1760.500 2917.600 1791.140 ;
        RECT 2.365 1758.500 2917.200 1760.500 ;
        RECT 2.365 1727.860 2917.600 1758.500 ;
        RECT 2.800 1725.860 2917.600 1727.860 ;
        RECT 2.365 1693.860 2917.600 1725.860 ;
        RECT 2.365 1691.860 2917.200 1693.860 ;
        RECT 2.365 1662.580 2917.600 1691.860 ;
        RECT 2.800 1660.580 2917.600 1662.580 ;
        RECT 2.365 1627.220 2917.600 1660.580 ;
        RECT 2.365 1625.220 2917.200 1627.220 ;
        RECT 2.365 1597.300 2917.600 1625.220 ;
        RECT 2.800 1595.300 2917.600 1597.300 ;
        RECT 2.365 1561.260 2917.600 1595.300 ;
        RECT 2.365 1559.260 2917.200 1561.260 ;
        RECT 2.365 1532.020 2917.600 1559.260 ;
        RECT 2.800 1530.020 2917.600 1532.020 ;
        RECT 2.365 1494.620 2917.600 1530.020 ;
        RECT 2.365 1492.620 2917.200 1494.620 ;
        RECT 2.365 1466.740 2917.600 1492.620 ;
        RECT 2.800 1464.740 2917.600 1466.740 ;
        RECT 2.365 1427.980 2917.600 1464.740 ;
        RECT 2.365 1425.980 2917.200 1427.980 ;
        RECT 2.365 1401.460 2917.600 1425.980 ;
        RECT 2.800 1399.460 2917.600 1401.460 ;
        RECT 2.365 1362.020 2917.600 1399.460 ;
        RECT 2.365 1360.020 2917.200 1362.020 ;
        RECT 2.365 1336.860 2917.600 1360.020 ;
        RECT 2.800 1334.860 2917.600 1336.860 ;
        RECT 2.365 1295.380 2917.600 1334.860 ;
        RECT 2.365 1293.380 2917.200 1295.380 ;
        RECT 2.365 1271.580 2917.600 1293.380 ;
        RECT 2.800 1269.580 2917.600 1271.580 ;
        RECT 2.365 1228.740 2917.600 1269.580 ;
        RECT 2.365 1226.740 2917.200 1228.740 ;
        RECT 2.365 1206.300 2917.600 1226.740 ;
        RECT 2.800 1204.300 2917.600 1206.300 ;
        RECT 2.365 1162.780 2917.600 1204.300 ;
        RECT 2.365 1160.780 2917.200 1162.780 ;
        RECT 2.365 1141.020 2917.600 1160.780 ;
        RECT 2.800 1139.020 2917.600 1141.020 ;
        RECT 2.365 1096.140 2917.600 1139.020 ;
        RECT 2.365 1094.140 2917.200 1096.140 ;
        RECT 2.365 1075.740 2917.600 1094.140 ;
        RECT 2.800 1073.740 2917.600 1075.740 ;
        RECT 2.365 1029.500 2917.600 1073.740 ;
        RECT 2.365 1027.500 2917.200 1029.500 ;
        RECT 2.365 1010.460 2917.600 1027.500 ;
        RECT 2.800 1008.460 2917.600 1010.460 ;
        RECT 2.365 963.540 2917.600 1008.460 ;
        RECT 2.365 961.540 2917.200 963.540 ;
        RECT 2.365 945.180 2917.600 961.540 ;
        RECT 2.800 943.180 2917.600 945.180 ;
        RECT 2.365 896.900 2917.600 943.180 ;
        RECT 2.365 894.900 2917.200 896.900 ;
        RECT 2.365 880.580 2917.600 894.900 ;
        RECT 2.800 878.580 2917.600 880.580 ;
        RECT 2.365 830.260 2917.600 878.580 ;
        RECT 2.365 828.260 2917.200 830.260 ;
        RECT 2.365 815.300 2917.600 828.260 ;
        RECT 2.800 813.300 2917.600 815.300 ;
        RECT 2.365 764.300 2917.600 813.300 ;
        RECT 2.365 762.300 2917.200 764.300 ;
        RECT 2.365 750.020 2917.600 762.300 ;
        RECT 2.800 748.020 2917.600 750.020 ;
        RECT 2.365 697.660 2917.600 748.020 ;
        RECT 2.365 695.660 2917.200 697.660 ;
        RECT 2.365 684.740 2917.600 695.660 ;
        RECT 2.800 682.740 2917.600 684.740 ;
        RECT 2.365 631.020 2917.600 682.740 ;
        RECT 2.365 629.020 2917.200 631.020 ;
        RECT 2.365 619.460 2917.600 629.020 ;
        RECT 2.800 617.460 2917.600 619.460 ;
        RECT 2.365 565.060 2917.600 617.460 ;
        RECT 2.365 563.060 2917.200 565.060 ;
        RECT 2.365 554.180 2917.600 563.060 ;
        RECT 2.800 552.180 2917.600 554.180 ;
        RECT 2.365 498.420 2917.600 552.180 ;
        RECT 2.365 496.420 2917.200 498.420 ;
        RECT 2.365 488.900 2917.600 496.420 ;
        RECT 2.800 486.900 2917.600 488.900 ;
        RECT 2.365 431.780 2917.600 486.900 ;
        RECT 2.365 429.780 2917.200 431.780 ;
        RECT 2.365 424.300 2917.600 429.780 ;
        RECT 2.800 422.300 2917.600 424.300 ;
        RECT 2.365 365.820 2917.600 422.300 ;
        RECT 2.365 363.820 2917.200 365.820 ;
        RECT 2.365 359.020 2917.600 363.820 ;
        RECT 2.800 357.020 2917.600 359.020 ;
        RECT 2.365 299.180 2917.600 357.020 ;
        RECT 2.365 297.180 2917.200 299.180 ;
        RECT 2.365 293.740 2917.600 297.180 ;
        RECT 2.800 291.740 2917.600 293.740 ;
        RECT 2.365 232.540 2917.600 291.740 ;
        RECT 2.365 230.540 2917.200 232.540 ;
        RECT 2.365 228.460 2917.600 230.540 ;
        RECT 2.800 226.460 2917.600 228.460 ;
        RECT 2.365 166.580 2917.600 226.460 ;
        RECT 2.365 164.580 2917.200 166.580 ;
        RECT 2.365 163.180 2917.600 164.580 ;
        RECT 2.800 161.180 2917.600 163.180 ;
        RECT 2.365 99.940 2917.600 161.180 ;
        RECT 2.365 97.940 2917.200 99.940 ;
        RECT 2.365 97.900 2917.600 97.940 ;
        RECT 2.800 95.900 2917.600 97.900 ;
        RECT 2.365 33.980 2917.600 95.900 ;
        RECT 2.365 33.300 2917.200 33.980 ;
        RECT 2.800 31.980 2917.200 33.300 ;
        RECT 2.800 31.300 2917.600 31.980 ;
        RECT 2.365 7.655 2917.600 31.300 ;
      LAYER met4 ;
        RECT 6.735 2203.280 8.570 3507.945 ;
        RECT 12.470 2203.520 27.170 3507.945 ;
        RECT 31.070 2203.520 45.770 3507.945 ;
        RECT 49.670 2203.520 64.370 3507.945 ;
        RECT 68.270 2203.520 98.570 3507.945 ;
        RECT 12.470 2203.280 98.570 2203.520 ;
        RECT 102.470 2203.520 117.170 3507.945 ;
        RECT 121.070 2203.520 135.770 3507.945 ;
        RECT 139.670 2203.520 154.370 3507.945 ;
        RECT 158.270 2203.520 188.570 3507.945 ;
        RECT 102.470 2203.280 188.570 2203.520 ;
        RECT 192.470 2203.520 207.170 3507.945 ;
        RECT 211.070 2203.520 225.770 3507.945 ;
        RECT 229.670 2203.520 244.370 3507.945 ;
        RECT 248.270 2203.520 278.570 3507.945 ;
        RECT 192.470 2203.280 278.570 2203.520 ;
        RECT 282.470 2203.520 297.170 3507.945 ;
        RECT 301.070 2203.520 315.770 3507.945 ;
        RECT 319.670 2203.520 334.370 3507.945 ;
        RECT 338.270 2203.520 368.570 3507.945 ;
        RECT 282.470 2203.280 368.570 2203.520 ;
        RECT 372.470 2203.520 387.170 3507.945 ;
        RECT 391.070 2203.520 405.770 3507.945 ;
        RECT 409.670 2203.520 424.370 3507.945 ;
        RECT 428.270 2203.520 458.570 3507.945 ;
        RECT 372.470 2203.280 458.570 2203.520 ;
        RECT 462.470 2203.520 477.170 3507.945 ;
        RECT 481.070 2203.520 495.770 3507.945 ;
        RECT 499.670 2203.520 514.370 3507.945 ;
        RECT 518.270 2203.520 548.570 3507.945 ;
        RECT 462.470 2203.280 548.570 2203.520 ;
        RECT 552.470 2203.520 567.170 3507.945 ;
        RECT 571.070 2203.520 585.770 3507.945 ;
        RECT 589.670 2203.520 604.370 3507.945 ;
        RECT 608.270 3488.240 638.570 3507.945 ;
        RECT 642.470 3488.480 657.170 3507.945 ;
        RECT 661.070 3488.480 675.770 3507.945 ;
        RECT 679.670 3488.480 694.370 3507.945 ;
        RECT 698.270 3488.480 728.570 3507.945 ;
        RECT 642.470 3488.240 728.570 3488.480 ;
        RECT 732.470 3488.480 747.170 3507.945 ;
        RECT 751.070 3488.480 765.770 3507.945 ;
        RECT 769.670 3488.480 784.370 3507.945 ;
        RECT 788.270 3488.480 818.570 3507.945 ;
        RECT 732.470 3488.240 818.570 3488.480 ;
        RECT 822.470 3488.480 837.170 3507.945 ;
        RECT 841.070 3488.480 855.770 3507.945 ;
        RECT 859.670 3488.480 874.370 3507.945 ;
        RECT 878.270 3488.480 908.570 3507.945 ;
        RECT 822.470 3488.240 908.570 3488.480 ;
        RECT 912.470 3488.480 927.170 3507.945 ;
        RECT 931.070 3488.480 945.770 3507.945 ;
        RECT 949.670 3488.480 964.370 3507.945 ;
        RECT 968.270 3488.480 998.570 3507.945 ;
        RECT 912.470 3488.240 998.570 3488.480 ;
        RECT 1002.470 3488.480 1017.170 3507.945 ;
        RECT 1021.070 3488.480 1035.770 3507.945 ;
        RECT 1039.670 3488.480 1054.370 3507.945 ;
        RECT 1058.270 3488.480 1088.570 3507.945 ;
        RECT 1002.470 3488.240 1088.570 3488.480 ;
        RECT 1092.470 3488.480 1107.170 3507.945 ;
        RECT 1111.070 3488.480 1125.770 3507.945 ;
        RECT 1129.670 3488.480 1144.370 3507.945 ;
        RECT 1148.270 3488.480 1178.570 3507.945 ;
        RECT 1092.470 3488.240 1178.570 3488.480 ;
        RECT 1182.470 3488.480 1197.170 3507.945 ;
        RECT 1201.070 3488.480 1215.770 3507.945 ;
        RECT 1219.670 3488.480 1234.370 3507.945 ;
        RECT 1238.270 3488.480 1268.570 3507.945 ;
        RECT 1182.470 3488.240 1268.570 3488.480 ;
        RECT 1272.470 3488.480 1287.170 3507.945 ;
        RECT 1291.070 3488.480 1305.770 3507.945 ;
        RECT 1309.670 3488.480 1324.370 3507.945 ;
        RECT 1328.270 3488.480 1358.570 3507.945 ;
        RECT 1272.470 3488.240 1358.570 3488.480 ;
        RECT 1362.470 3488.480 1377.170 3507.945 ;
        RECT 1381.070 3488.480 1395.770 3507.945 ;
        RECT 1399.670 3488.480 1414.370 3507.945 ;
        RECT 1418.270 3488.480 1448.570 3507.945 ;
        RECT 1362.470 3488.240 1448.570 3488.480 ;
        RECT 1452.470 3488.480 1467.170 3507.945 ;
        RECT 1471.070 3488.480 1485.770 3507.945 ;
        RECT 1489.670 3488.480 1504.370 3507.945 ;
        RECT 1508.270 3488.480 1538.570 3507.945 ;
        RECT 1452.470 3488.240 1538.570 3488.480 ;
        RECT 1542.470 3488.480 1557.170 3507.945 ;
        RECT 1561.070 3488.480 1575.770 3507.945 ;
        RECT 1579.670 3488.480 1594.370 3507.945 ;
        RECT 1598.270 3488.480 1628.570 3507.945 ;
        RECT 1542.470 3488.240 1628.570 3488.480 ;
        RECT 1632.470 3488.480 1647.170 3507.945 ;
        RECT 1651.070 3488.480 1665.770 3507.945 ;
        RECT 1669.670 3488.480 1684.370 3507.945 ;
        RECT 1688.270 3488.480 1718.570 3507.945 ;
        RECT 1632.470 3488.240 1718.570 3488.480 ;
        RECT 1722.470 3488.480 1737.170 3507.945 ;
        RECT 1741.070 3488.480 1755.770 3507.945 ;
        RECT 1759.670 3488.480 1774.370 3507.945 ;
        RECT 1778.270 3488.480 1808.570 3507.945 ;
        RECT 1722.470 3488.240 1808.570 3488.480 ;
        RECT 1812.470 3488.480 1827.170 3507.945 ;
        RECT 1831.070 3488.480 1845.770 3507.945 ;
        RECT 1849.670 3488.480 1864.370 3507.945 ;
        RECT 1868.270 3488.480 1898.570 3507.945 ;
        RECT 1812.470 3488.240 1898.570 3488.480 ;
        RECT 1902.470 3488.480 1917.170 3507.945 ;
        RECT 1921.070 3488.480 1935.770 3507.945 ;
        RECT 1939.670 3488.480 1954.370 3507.945 ;
        RECT 1958.270 3488.480 1988.570 3507.945 ;
        RECT 1902.470 3488.240 1988.570 3488.480 ;
        RECT 1992.470 3488.480 2007.170 3507.945 ;
        RECT 2011.070 3488.480 2025.770 3507.945 ;
        RECT 2029.670 3488.480 2044.370 3507.945 ;
        RECT 2048.270 3488.480 2078.570 3507.945 ;
        RECT 1992.470 3488.240 2078.570 3488.480 ;
        RECT 2082.470 3488.480 2097.170 3507.945 ;
        RECT 2101.070 3488.480 2115.770 3507.945 ;
        RECT 2119.670 3488.480 2134.370 3507.945 ;
        RECT 2138.270 3488.480 2168.570 3507.945 ;
        RECT 2082.470 3488.240 2168.570 3488.480 ;
        RECT 2172.470 3488.480 2187.170 3507.945 ;
        RECT 2191.070 3488.480 2205.770 3507.945 ;
        RECT 2209.670 3488.480 2224.370 3507.945 ;
        RECT 2228.270 3488.480 2258.570 3507.945 ;
        RECT 2172.470 3488.240 2258.570 3488.480 ;
        RECT 2262.470 3488.480 2277.170 3507.945 ;
        RECT 2281.070 3488.480 2295.770 3507.945 ;
        RECT 2262.470 3488.240 2295.770 3488.480 ;
        RECT 608.270 2482.160 2295.770 3488.240 ;
        RECT 608.270 2203.520 638.570 2482.160 ;
        RECT 552.470 2203.280 638.570 2203.520 ;
        RECT 642.470 2481.920 728.570 2482.160 ;
        RECT 642.470 2203.520 657.170 2481.920 ;
        RECT 661.070 2203.520 675.770 2481.920 ;
        RECT 679.670 2203.520 694.370 2481.920 ;
        RECT 642.470 2203.280 694.370 2203.520 ;
        RECT 6.735 1584.560 694.370 2203.280 ;
        RECT 6.735 1137.040 8.570 1584.560 ;
        RECT 12.470 1584.320 98.570 1584.560 ;
        RECT 12.470 1137.280 27.170 1584.320 ;
        RECT 31.070 1137.280 45.770 1584.320 ;
        RECT 49.670 1137.280 64.370 1584.320 ;
        RECT 68.270 1137.280 98.570 1584.320 ;
        RECT 12.470 1137.040 98.570 1137.280 ;
        RECT 102.470 1584.320 188.570 1584.560 ;
        RECT 102.470 1137.280 117.170 1584.320 ;
        RECT 121.070 1137.280 135.770 1584.320 ;
        RECT 139.670 1137.280 154.370 1584.320 ;
        RECT 158.270 1137.280 188.570 1584.320 ;
        RECT 102.470 1137.040 188.570 1137.280 ;
        RECT 192.470 1584.320 278.570 1584.560 ;
        RECT 192.470 1137.280 207.170 1584.320 ;
        RECT 211.070 1137.280 225.770 1584.320 ;
        RECT 229.670 1137.280 244.370 1584.320 ;
        RECT 248.270 1137.280 278.570 1584.320 ;
        RECT 192.470 1137.040 278.570 1137.280 ;
        RECT 282.470 1584.320 368.570 1584.560 ;
        RECT 282.470 1137.280 297.170 1584.320 ;
        RECT 301.070 1137.280 315.770 1584.320 ;
        RECT 319.670 1137.280 334.370 1584.320 ;
        RECT 338.270 1137.280 368.570 1584.320 ;
        RECT 282.470 1137.040 368.570 1137.280 ;
        RECT 372.470 1584.320 458.570 1584.560 ;
        RECT 372.470 1137.280 387.170 1584.320 ;
        RECT 391.070 1137.280 405.770 1584.320 ;
        RECT 409.670 1137.280 424.370 1584.320 ;
        RECT 428.270 1137.280 458.570 1584.320 ;
        RECT 372.470 1137.040 458.570 1137.280 ;
        RECT 462.470 1584.320 548.570 1584.560 ;
        RECT 462.470 1137.280 477.170 1584.320 ;
        RECT 481.070 1137.280 495.770 1584.320 ;
        RECT 499.670 1137.280 514.370 1584.320 ;
        RECT 518.270 1137.280 548.570 1584.320 ;
        RECT 462.470 1137.040 548.570 1137.280 ;
        RECT 552.470 1584.320 638.570 1584.560 ;
        RECT 552.470 1137.280 567.170 1584.320 ;
        RECT 571.070 1137.280 585.770 1584.320 ;
        RECT 589.670 1137.280 604.370 1584.320 ;
        RECT 608.270 1137.280 638.570 1584.320 ;
        RECT 552.470 1137.040 638.570 1137.280 ;
        RECT 642.470 1584.320 694.370 1584.560 ;
        RECT 642.470 1137.280 657.170 1584.320 ;
        RECT 661.070 1137.280 675.770 1584.320 ;
        RECT 679.670 1137.280 694.370 1584.320 ;
        RECT 642.470 1137.040 694.370 1137.280 ;
        RECT 6.735 518.320 694.370 1137.040 ;
        RECT 6.735 235.600 8.570 518.320 ;
        RECT 12.470 518.080 98.570 518.320 ;
        RECT 12.470 235.840 27.170 518.080 ;
        RECT 31.070 235.840 45.770 518.080 ;
        RECT 49.670 235.840 64.370 518.080 ;
        RECT 68.270 235.840 98.570 518.080 ;
        RECT 12.470 235.600 98.570 235.840 ;
        RECT 102.470 518.080 188.570 518.320 ;
        RECT 102.470 235.840 117.170 518.080 ;
        RECT 121.070 235.840 135.770 518.080 ;
        RECT 139.670 235.840 154.370 518.080 ;
        RECT 158.270 235.840 188.570 518.080 ;
        RECT 102.470 235.600 188.570 235.840 ;
        RECT 192.470 518.080 278.570 518.320 ;
        RECT 192.470 235.840 207.170 518.080 ;
        RECT 211.070 235.840 225.770 518.080 ;
        RECT 229.670 235.840 244.370 518.080 ;
        RECT 248.270 235.840 278.570 518.080 ;
        RECT 192.470 235.600 278.570 235.840 ;
        RECT 282.470 518.080 368.570 518.320 ;
        RECT 282.470 235.840 297.170 518.080 ;
        RECT 301.070 235.840 315.770 518.080 ;
        RECT 319.670 235.840 334.370 518.080 ;
        RECT 338.270 235.840 368.570 518.080 ;
        RECT 282.470 235.600 368.570 235.840 ;
        RECT 372.470 518.080 458.570 518.320 ;
        RECT 372.470 235.840 387.170 518.080 ;
        RECT 391.070 235.840 405.770 518.080 ;
        RECT 409.670 235.840 424.370 518.080 ;
        RECT 428.270 235.840 458.570 518.080 ;
        RECT 372.470 235.600 458.570 235.840 ;
        RECT 462.470 518.080 548.570 518.320 ;
        RECT 462.470 235.840 477.170 518.080 ;
        RECT 481.070 235.840 495.770 518.080 ;
        RECT 499.670 235.840 514.370 518.080 ;
        RECT 518.270 235.840 548.570 518.080 ;
        RECT 462.470 235.600 548.570 235.840 ;
        RECT 552.470 518.080 638.570 518.320 ;
        RECT 552.470 235.840 567.170 518.080 ;
        RECT 571.070 235.840 585.770 518.080 ;
        RECT 589.670 235.840 604.370 518.080 ;
        RECT 608.270 235.840 638.570 518.080 ;
        RECT 552.470 235.600 638.570 235.840 ;
        RECT 642.470 518.080 694.370 518.320 ;
        RECT 642.470 235.840 657.170 518.080 ;
        RECT 661.070 235.840 675.770 518.080 ;
        RECT 679.670 235.840 694.370 518.080 ;
        RECT 698.270 235.840 728.570 2481.920 ;
        RECT 642.470 235.600 728.570 235.840 ;
        RECT 732.470 2481.920 818.570 2482.160 ;
        RECT 732.470 235.840 747.170 2481.920 ;
        RECT 751.070 235.840 765.770 2481.920 ;
        RECT 769.670 235.840 784.370 2481.920 ;
        RECT 788.270 235.840 818.570 2481.920 ;
        RECT 732.470 235.600 818.570 235.840 ;
        RECT 822.470 2481.920 908.570 2482.160 ;
        RECT 822.470 235.840 837.170 2481.920 ;
        RECT 841.070 235.840 855.770 2481.920 ;
        RECT 859.670 235.840 874.370 2481.920 ;
        RECT 878.270 235.840 908.570 2481.920 ;
        RECT 822.470 235.600 908.570 235.840 ;
        RECT 912.470 2481.920 998.570 2482.160 ;
        RECT 912.470 235.840 927.170 2481.920 ;
        RECT 931.070 235.840 945.770 2481.920 ;
        RECT 949.670 235.840 964.370 2481.920 ;
        RECT 968.270 235.840 998.570 2481.920 ;
        RECT 912.470 235.600 998.570 235.840 ;
        RECT 1002.470 2481.920 1088.570 2482.160 ;
        RECT 1002.470 235.840 1017.170 2481.920 ;
        RECT 1021.070 235.840 1035.770 2481.920 ;
        RECT 1039.670 235.840 1054.370 2481.920 ;
        RECT 1058.270 235.840 1088.570 2481.920 ;
        RECT 1002.470 235.600 1088.570 235.840 ;
        RECT 1092.470 2481.920 1178.570 2482.160 ;
        RECT 1092.470 235.840 1107.170 2481.920 ;
        RECT 1111.070 235.840 1125.770 2481.920 ;
        RECT 1129.670 235.840 1144.370 2481.920 ;
        RECT 1148.270 235.840 1178.570 2481.920 ;
        RECT 1092.470 235.600 1178.570 235.840 ;
        RECT 1182.470 2481.920 1268.570 2482.160 ;
        RECT 1182.470 235.840 1197.170 2481.920 ;
        RECT 1201.070 235.840 1215.770 2481.920 ;
        RECT 1219.670 235.840 1234.370 2481.920 ;
        RECT 1238.270 235.840 1268.570 2481.920 ;
        RECT 1182.470 235.600 1268.570 235.840 ;
        RECT 6.735 31.440 1268.570 235.600 ;
        RECT 6.735 7.655 8.570 31.440 ;
        RECT 12.470 31.200 98.570 31.440 ;
        RECT 12.470 7.655 27.170 31.200 ;
        RECT 31.070 7.655 45.770 31.200 ;
        RECT 49.670 7.655 64.370 31.200 ;
        RECT 68.270 7.655 98.570 31.200 ;
        RECT 102.470 31.200 188.570 31.440 ;
        RECT 102.470 7.655 117.170 31.200 ;
        RECT 121.070 7.655 135.770 31.200 ;
        RECT 139.670 7.655 154.370 31.200 ;
        RECT 158.270 7.655 188.570 31.200 ;
        RECT 192.470 31.200 278.570 31.440 ;
        RECT 192.470 7.655 207.170 31.200 ;
        RECT 211.070 7.655 225.770 31.200 ;
        RECT 229.670 7.655 244.370 31.200 ;
        RECT 248.270 7.655 278.570 31.200 ;
        RECT 282.470 31.200 368.570 31.440 ;
        RECT 282.470 7.655 297.170 31.200 ;
        RECT 301.070 7.655 315.770 31.200 ;
        RECT 319.670 7.655 334.370 31.200 ;
        RECT 338.270 7.655 368.570 31.200 ;
        RECT 372.470 31.200 458.570 31.440 ;
        RECT 372.470 7.655 387.170 31.200 ;
        RECT 391.070 7.655 405.770 31.200 ;
        RECT 409.670 7.655 424.370 31.200 ;
        RECT 428.270 7.655 458.570 31.200 ;
        RECT 462.470 31.200 548.570 31.440 ;
        RECT 462.470 7.655 477.170 31.200 ;
        RECT 481.070 7.655 495.770 31.200 ;
        RECT 499.670 7.655 514.370 31.200 ;
        RECT 518.270 7.655 548.570 31.200 ;
        RECT 552.470 31.200 638.570 31.440 ;
        RECT 552.470 7.655 567.170 31.200 ;
        RECT 571.070 7.655 585.770 31.200 ;
        RECT 589.670 7.655 604.370 31.200 ;
        RECT 608.270 7.655 638.570 31.200 ;
        RECT 642.470 31.200 728.570 31.440 ;
        RECT 642.470 7.655 657.170 31.200 ;
        RECT 661.070 7.655 675.770 31.200 ;
        RECT 679.670 7.655 694.370 31.200 ;
        RECT 698.270 7.655 728.570 31.200 ;
        RECT 732.470 31.200 818.570 31.440 ;
        RECT 732.470 7.655 747.170 31.200 ;
        RECT 751.070 7.655 765.770 31.200 ;
        RECT 769.670 7.655 784.370 31.200 ;
        RECT 788.270 7.655 818.570 31.200 ;
        RECT 822.470 31.200 908.570 31.440 ;
        RECT 822.470 7.655 837.170 31.200 ;
        RECT 841.070 7.655 855.770 31.200 ;
        RECT 859.670 7.655 874.370 31.200 ;
        RECT 878.270 7.655 908.570 31.200 ;
        RECT 912.470 31.200 998.570 31.440 ;
        RECT 912.470 7.655 927.170 31.200 ;
        RECT 931.070 7.655 945.770 31.200 ;
        RECT 949.670 7.655 964.370 31.200 ;
        RECT 968.270 7.655 998.570 31.200 ;
        RECT 1002.470 31.200 1088.570 31.440 ;
        RECT 1002.470 7.655 1017.170 31.200 ;
        RECT 1021.070 7.655 1035.770 31.200 ;
        RECT 1039.670 7.655 1054.370 31.200 ;
        RECT 1058.270 7.655 1088.570 31.200 ;
        RECT 1092.470 31.200 1178.570 31.440 ;
        RECT 1092.470 7.655 1107.170 31.200 ;
        RECT 1111.070 7.655 1125.770 31.200 ;
        RECT 1129.670 7.655 1144.370 31.200 ;
        RECT 1148.270 7.655 1178.570 31.200 ;
        RECT 1182.470 31.200 1268.570 31.440 ;
        RECT 1182.470 7.655 1197.170 31.200 ;
        RECT 1201.070 7.655 1215.770 31.200 ;
        RECT 1219.670 7.655 1234.370 31.200 ;
        RECT 1238.270 7.655 1268.570 31.200 ;
        RECT 1272.470 2481.920 1358.570 2482.160 ;
        RECT 1272.470 7.655 1287.170 2481.920 ;
        RECT 1291.070 7.655 1305.770 2481.920 ;
        RECT 1309.670 7.655 1324.370 2481.920 ;
        RECT 1328.270 7.655 1358.570 2481.920 ;
        RECT 1362.470 2481.920 1448.570 2482.160 ;
        RECT 1362.470 7.655 1377.170 2481.920 ;
        RECT 1381.070 7.655 1395.770 2481.920 ;
        RECT 1399.670 7.655 1414.370 2481.920 ;
        RECT 1418.270 7.655 1448.570 2481.920 ;
        RECT 1452.470 2481.920 1538.570 2482.160 ;
        RECT 1452.470 7.655 1467.170 2481.920 ;
        RECT 1471.070 7.655 1485.770 2481.920 ;
        RECT 1489.670 7.655 1504.370 2481.920 ;
        RECT 1508.270 7.655 1538.570 2481.920 ;
        RECT 1542.470 2481.920 1628.570 2482.160 ;
        RECT 1542.470 7.655 1557.170 2481.920 ;
        RECT 1561.070 7.655 1575.770 2481.920 ;
        RECT 1579.670 7.655 1594.370 2481.920 ;
        RECT 1598.270 7.655 1628.570 2481.920 ;
        RECT 1632.470 2481.920 1718.570 2482.160 ;
        RECT 1632.470 7.655 1647.170 2481.920 ;
        RECT 1651.070 235.840 1665.770 2481.920 ;
        RECT 1669.670 235.840 1684.370 2481.920 ;
        RECT 1688.270 1945.440 1718.570 2481.920 ;
        RECT 1722.470 2481.920 1808.570 2482.160 ;
        RECT 1722.470 1945.680 1737.170 2481.920 ;
        RECT 1741.070 1945.680 1755.770 2481.920 ;
        RECT 1759.670 1945.680 1774.370 2481.920 ;
        RECT 1778.270 1945.680 1808.570 2481.920 ;
        RECT 1722.470 1945.440 1808.570 1945.680 ;
        RECT 1812.470 2481.920 1898.570 2482.160 ;
        RECT 1812.470 1945.680 1827.170 2481.920 ;
        RECT 1831.070 1945.680 1845.770 2481.920 ;
        RECT 1849.670 1945.680 1864.370 2481.920 ;
        RECT 1868.270 1945.680 1898.570 2481.920 ;
        RECT 1812.470 1945.440 1898.570 1945.680 ;
        RECT 1902.470 2481.920 1988.570 2482.160 ;
        RECT 1902.470 1945.680 1917.170 2481.920 ;
        RECT 1921.070 1945.680 1935.770 2481.920 ;
        RECT 1939.670 1945.680 1954.370 2481.920 ;
        RECT 1958.270 1945.680 1988.570 2481.920 ;
        RECT 1902.470 1945.440 1988.570 1945.680 ;
        RECT 1992.470 2481.920 2078.570 2482.160 ;
        RECT 1992.470 1945.680 2007.170 2481.920 ;
        RECT 2011.070 1945.680 2025.770 2481.920 ;
        RECT 2029.670 1945.680 2044.370 2481.920 ;
        RECT 2048.270 1945.680 2078.570 2481.920 ;
        RECT 1992.470 1945.440 2078.570 1945.680 ;
        RECT 2082.470 2481.920 2168.570 2482.160 ;
        RECT 2082.470 1945.680 2097.170 2481.920 ;
        RECT 2101.070 1945.680 2115.770 2481.920 ;
        RECT 2119.670 1945.680 2134.370 2481.920 ;
        RECT 2138.270 1945.680 2168.570 2481.920 ;
        RECT 2082.470 1945.440 2168.570 1945.680 ;
        RECT 2172.470 2481.920 2258.570 2482.160 ;
        RECT 2172.470 1945.680 2187.170 2481.920 ;
        RECT 2191.070 1945.680 2205.770 2481.920 ;
        RECT 2209.670 1945.680 2224.370 2481.920 ;
        RECT 2228.270 1945.680 2258.570 2481.920 ;
        RECT 2172.470 1945.440 2258.570 1945.680 ;
        RECT 2262.470 2481.920 2295.770 2482.160 ;
        RECT 2262.470 1945.680 2277.170 2481.920 ;
        RECT 2281.070 1945.680 2295.770 2481.920 ;
        RECT 2299.670 1945.680 2314.370 3507.945 ;
        RECT 2318.270 1945.680 2348.570 3507.945 ;
        RECT 2262.470 1945.440 2348.570 1945.680 ;
        RECT 2352.470 1945.680 2367.170 3507.945 ;
        RECT 2371.070 1945.680 2385.770 3507.945 ;
        RECT 2389.670 1945.680 2404.370 3507.945 ;
        RECT 2408.270 1945.680 2438.570 3507.945 ;
        RECT 2352.470 1945.440 2438.570 1945.680 ;
        RECT 2442.470 1945.680 2457.170 3507.945 ;
        RECT 2461.070 1945.680 2475.770 3507.945 ;
        RECT 2479.670 1945.680 2494.370 3507.945 ;
        RECT 2498.270 1945.680 2528.570 3507.945 ;
        RECT 2442.470 1945.440 2528.570 1945.680 ;
        RECT 2532.470 1945.680 2547.170 3507.945 ;
        RECT 2551.070 1945.680 2565.770 3507.945 ;
        RECT 2569.670 1945.680 2584.370 3507.945 ;
        RECT 2588.270 1945.680 2618.570 3507.945 ;
        RECT 2532.470 1945.440 2618.570 1945.680 ;
        RECT 2622.470 1945.680 2637.170 3507.945 ;
        RECT 2641.070 1945.680 2655.770 3507.945 ;
        RECT 2659.670 1945.680 2674.370 3507.945 ;
        RECT 2678.270 1945.680 2708.570 3507.945 ;
        RECT 2622.470 1945.440 2708.570 1945.680 ;
        RECT 2712.470 1945.680 2727.170 3507.945 ;
        RECT 2731.070 1945.680 2745.770 3507.945 ;
        RECT 2749.670 1945.680 2764.370 3507.945 ;
        RECT 2768.270 1945.680 2798.570 3507.945 ;
        RECT 2712.470 1945.440 2798.570 1945.680 ;
        RECT 2802.470 1945.680 2817.170 3507.945 ;
        RECT 2821.070 1945.680 2835.770 3507.945 ;
        RECT 2839.670 1945.680 2848.025 3507.945 ;
        RECT 2802.470 1945.440 2848.025 1945.680 ;
        RECT 1688.270 776.720 2848.025 1945.440 ;
        RECT 1688.270 235.840 1718.570 776.720 ;
        RECT 1651.070 235.600 1718.570 235.840 ;
        RECT 1722.470 776.480 1808.570 776.720 ;
        RECT 1722.470 235.840 1737.170 776.480 ;
        RECT 1741.070 235.840 1755.770 776.480 ;
        RECT 1759.670 235.840 1774.370 776.480 ;
        RECT 1778.270 235.840 1808.570 776.480 ;
        RECT 1722.470 235.600 1808.570 235.840 ;
        RECT 1812.470 776.480 1898.570 776.720 ;
        RECT 1812.470 235.840 1827.170 776.480 ;
        RECT 1831.070 235.840 1845.770 776.480 ;
        RECT 1849.670 235.840 1864.370 776.480 ;
        RECT 1868.270 235.840 1898.570 776.480 ;
        RECT 1812.470 235.600 1898.570 235.840 ;
        RECT 1902.470 776.480 1988.570 776.720 ;
        RECT 1902.470 235.840 1917.170 776.480 ;
        RECT 1921.070 235.840 1935.770 776.480 ;
        RECT 1939.670 235.840 1954.370 776.480 ;
        RECT 1958.270 235.840 1988.570 776.480 ;
        RECT 1902.470 235.600 1988.570 235.840 ;
        RECT 1992.470 776.480 2078.570 776.720 ;
        RECT 1992.470 235.840 2007.170 776.480 ;
        RECT 2011.070 235.840 2025.770 776.480 ;
        RECT 2029.670 235.840 2044.370 776.480 ;
        RECT 2048.270 235.840 2078.570 776.480 ;
        RECT 1992.470 235.600 2078.570 235.840 ;
        RECT 2082.470 776.480 2168.570 776.720 ;
        RECT 2082.470 235.840 2097.170 776.480 ;
        RECT 2101.070 235.840 2115.770 776.480 ;
        RECT 2119.670 235.840 2134.370 776.480 ;
        RECT 2138.270 235.840 2168.570 776.480 ;
        RECT 2082.470 235.600 2168.570 235.840 ;
        RECT 2172.470 776.480 2258.570 776.720 ;
        RECT 2172.470 235.840 2187.170 776.480 ;
        RECT 2191.070 235.840 2205.770 776.480 ;
        RECT 2209.670 235.840 2224.370 776.480 ;
        RECT 2228.270 235.840 2258.570 776.480 ;
        RECT 2172.470 235.600 2258.570 235.840 ;
        RECT 2262.470 776.480 2348.570 776.720 ;
        RECT 2262.470 235.840 2277.170 776.480 ;
        RECT 2281.070 235.840 2295.770 776.480 ;
        RECT 2299.670 235.840 2314.370 776.480 ;
        RECT 2318.270 235.840 2348.570 776.480 ;
        RECT 2262.470 235.600 2348.570 235.840 ;
        RECT 2352.470 776.480 2438.570 776.720 ;
        RECT 2352.470 235.840 2367.170 776.480 ;
        RECT 2371.070 235.840 2385.770 776.480 ;
        RECT 2389.670 235.840 2404.370 776.480 ;
        RECT 2408.270 235.840 2438.570 776.480 ;
        RECT 2352.470 235.600 2438.570 235.840 ;
        RECT 2442.470 776.480 2528.570 776.720 ;
        RECT 2442.470 235.840 2457.170 776.480 ;
        RECT 2461.070 235.840 2475.770 776.480 ;
        RECT 2479.670 235.840 2494.370 776.480 ;
        RECT 2498.270 235.840 2528.570 776.480 ;
        RECT 2442.470 235.600 2528.570 235.840 ;
        RECT 2532.470 776.480 2618.570 776.720 ;
        RECT 2532.470 235.840 2547.170 776.480 ;
        RECT 2551.070 235.840 2565.770 776.480 ;
        RECT 2569.670 235.840 2584.370 776.480 ;
        RECT 2588.270 235.840 2618.570 776.480 ;
        RECT 2532.470 235.600 2618.570 235.840 ;
        RECT 2622.470 776.480 2708.570 776.720 ;
        RECT 2622.470 235.840 2637.170 776.480 ;
        RECT 2641.070 235.840 2655.770 776.480 ;
        RECT 2659.670 235.840 2674.370 776.480 ;
        RECT 2678.270 235.840 2708.570 776.480 ;
        RECT 2622.470 235.600 2708.570 235.840 ;
        RECT 2712.470 776.480 2798.570 776.720 ;
        RECT 2712.470 235.840 2727.170 776.480 ;
        RECT 2731.070 235.840 2745.770 776.480 ;
        RECT 2749.670 235.840 2764.370 776.480 ;
        RECT 2768.270 235.840 2798.570 776.480 ;
        RECT 2712.470 235.600 2798.570 235.840 ;
        RECT 2802.470 776.480 2848.025 776.720 ;
        RECT 2802.470 235.840 2817.170 776.480 ;
        RECT 2821.070 235.840 2835.770 776.480 ;
        RECT 2839.670 235.840 2848.025 776.480 ;
        RECT 2802.470 235.600 2848.025 235.840 ;
        RECT 1651.070 31.440 2848.025 235.600 ;
        RECT 1651.070 31.200 1718.570 31.440 ;
        RECT 1651.070 7.655 1665.770 31.200 ;
        RECT 1669.670 7.655 1684.370 31.200 ;
        RECT 1688.270 7.655 1718.570 31.200 ;
        RECT 1722.470 31.200 1808.570 31.440 ;
        RECT 1722.470 7.655 1737.170 31.200 ;
        RECT 1741.070 7.655 1755.770 31.200 ;
        RECT 1759.670 7.655 1774.370 31.200 ;
        RECT 1778.270 7.655 1808.570 31.200 ;
        RECT 1812.470 31.200 1898.570 31.440 ;
        RECT 1812.470 7.655 1827.170 31.200 ;
        RECT 1831.070 7.655 1845.770 31.200 ;
        RECT 1849.670 7.655 1864.370 31.200 ;
        RECT 1868.270 7.655 1898.570 31.200 ;
        RECT 1902.470 31.200 1988.570 31.440 ;
        RECT 1902.470 7.655 1917.170 31.200 ;
        RECT 1921.070 7.655 1935.770 31.200 ;
        RECT 1939.670 7.655 1954.370 31.200 ;
        RECT 1958.270 7.655 1988.570 31.200 ;
        RECT 1992.470 31.200 2078.570 31.440 ;
        RECT 1992.470 7.655 2007.170 31.200 ;
        RECT 2011.070 7.655 2025.770 31.200 ;
        RECT 2029.670 7.655 2044.370 31.200 ;
        RECT 2048.270 7.655 2078.570 31.200 ;
        RECT 2082.470 31.200 2168.570 31.440 ;
        RECT 2082.470 7.655 2097.170 31.200 ;
        RECT 2101.070 7.655 2115.770 31.200 ;
        RECT 2119.670 7.655 2134.370 31.200 ;
        RECT 2138.270 7.655 2168.570 31.200 ;
        RECT 2172.470 31.200 2258.570 31.440 ;
        RECT 2172.470 7.655 2187.170 31.200 ;
        RECT 2191.070 7.655 2205.770 31.200 ;
        RECT 2209.670 7.655 2224.370 31.200 ;
        RECT 2228.270 7.655 2258.570 31.200 ;
        RECT 2262.470 31.200 2348.570 31.440 ;
        RECT 2262.470 7.655 2277.170 31.200 ;
        RECT 2281.070 7.655 2295.770 31.200 ;
        RECT 2299.670 7.655 2314.370 31.200 ;
        RECT 2318.270 7.655 2348.570 31.200 ;
        RECT 2352.470 31.200 2438.570 31.440 ;
        RECT 2352.470 7.655 2367.170 31.200 ;
        RECT 2371.070 7.655 2385.770 31.200 ;
        RECT 2389.670 7.655 2404.370 31.200 ;
        RECT 2408.270 7.655 2438.570 31.200 ;
        RECT 2442.470 31.200 2528.570 31.440 ;
        RECT 2442.470 7.655 2457.170 31.200 ;
        RECT 2461.070 7.655 2475.770 31.200 ;
        RECT 2479.670 7.655 2494.370 31.200 ;
        RECT 2498.270 7.655 2528.570 31.200 ;
        RECT 2532.470 31.200 2618.570 31.440 ;
        RECT 2532.470 7.655 2547.170 31.200 ;
        RECT 2551.070 7.655 2565.770 31.200 ;
        RECT 2569.670 7.655 2584.370 31.200 ;
        RECT 2588.270 7.655 2618.570 31.200 ;
        RECT 2622.470 31.200 2708.570 31.440 ;
        RECT 2622.470 7.655 2637.170 31.200 ;
        RECT 2641.070 7.655 2655.770 31.200 ;
        RECT 2659.670 7.655 2674.370 31.200 ;
        RECT 2678.270 7.655 2708.570 31.200 ;
        RECT 2712.470 31.200 2798.570 31.440 ;
        RECT 2712.470 7.655 2727.170 31.200 ;
        RECT 2731.070 7.655 2745.770 31.200 ;
        RECT 2749.670 7.655 2764.370 31.200 ;
        RECT 2768.270 7.655 2798.570 31.200 ;
        RECT 2802.470 31.200 2848.025 31.440 ;
        RECT 2802.470 7.655 2817.170 31.200 ;
        RECT 2821.070 7.655 2835.770 31.200 ;
        RECT 2839.670 7.655 2848.025 31.200 ;
      LAYER met5 ;
        RECT 14.380 3404.830 2781.500 3409.300 ;
        RECT 14.380 3386.230 2781.500 3398.530 ;
        RECT 14.380 3367.630 2781.500 3379.930 ;
        RECT 14.380 3348.790 2781.500 3361.330 ;
        RECT 14.380 3314.830 2781.500 3342.490 ;
        RECT 14.380 3296.230 2781.500 3308.530 ;
        RECT 14.380 3277.630 2781.500 3289.930 ;
        RECT 14.380 3258.790 2781.500 3271.330 ;
        RECT 14.380 3224.830 2781.500 3252.490 ;
        RECT 14.380 3206.230 2781.500 3218.530 ;
        RECT 14.380 3187.630 2781.500 3199.930 ;
        RECT 14.380 3168.790 2781.500 3181.330 ;
        RECT 14.380 3134.830 2781.500 3162.490 ;
        RECT 14.380 3116.230 2781.500 3128.530 ;
        RECT 14.380 3097.630 2781.500 3109.930 ;
        RECT 14.380 3078.790 2781.500 3091.330 ;
        RECT 14.380 3044.830 2781.500 3072.490 ;
        RECT 14.380 3026.230 2781.500 3038.530 ;
        RECT 14.380 3007.630 2781.500 3019.930 ;
        RECT 14.380 2988.790 2781.500 3001.330 ;
        RECT 14.380 2954.830 2781.500 2982.490 ;
        RECT 14.380 2936.230 2781.500 2948.530 ;
        RECT 14.380 2917.630 2781.500 2929.930 ;
        RECT 14.380 2898.790 2781.500 2911.330 ;
        RECT 14.380 2864.830 2781.500 2892.490 ;
        RECT 14.380 2846.230 2781.500 2858.530 ;
        RECT 14.380 2827.630 2781.500 2839.930 ;
        RECT 14.380 2808.790 2781.500 2821.330 ;
        RECT 14.380 2774.830 2781.500 2802.490 ;
        RECT 14.380 2756.230 2781.500 2768.530 ;
        RECT 14.380 2737.630 2781.500 2749.930 ;
        RECT 14.380 2718.790 2781.500 2731.330 ;
        RECT 14.380 2684.830 2781.500 2712.490 ;
        RECT 14.380 2666.230 2781.500 2678.530 ;
        RECT 14.380 2647.630 2781.500 2659.930 ;
        RECT 14.380 2628.790 2781.500 2641.330 ;
        RECT 14.380 2594.830 2781.500 2622.490 ;
        RECT 14.380 2576.230 2781.500 2588.530 ;
        RECT 14.380 2557.630 2781.500 2569.930 ;
        RECT 14.380 2538.790 2781.500 2551.330 ;
        RECT 14.380 2504.830 2781.500 2532.490 ;
        RECT 14.380 2486.230 2781.500 2498.530 ;
        RECT 14.380 2467.630 2781.500 2479.930 ;
        RECT 14.380 2448.790 2781.500 2461.330 ;
        RECT 14.380 2414.830 2781.500 2442.490 ;
        RECT 14.380 2396.230 2781.500 2408.530 ;
        RECT 14.380 2377.630 2781.500 2389.930 ;
        RECT 14.380 2358.790 2781.500 2371.330 ;
        RECT 14.380 2324.830 2781.500 2352.490 ;
        RECT 14.380 2306.230 2781.500 2318.530 ;
        RECT 14.380 2287.630 2781.500 2299.930 ;
        RECT 14.380 2268.790 2781.500 2281.330 ;
        RECT 14.380 2234.830 2781.500 2262.490 ;
        RECT 14.380 2216.230 2781.500 2228.530 ;
        RECT 14.380 2197.630 2781.500 2209.930 ;
        RECT 14.380 2178.790 2781.500 2191.330 ;
        RECT 14.380 2144.830 2781.500 2172.490 ;
        RECT 14.380 2126.230 2781.500 2138.530 ;
        RECT 14.380 2107.630 2781.500 2119.930 ;
        RECT 14.380 2088.790 2781.500 2101.330 ;
        RECT 14.380 2054.830 2781.500 2082.490 ;
        RECT 14.380 2036.230 2781.500 2048.530 ;
        RECT 14.380 2017.630 2781.500 2029.930 ;
        RECT 14.380 1998.790 2781.500 2011.330 ;
        RECT 14.380 1964.830 2781.500 1992.490 ;
        RECT 14.380 1946.230 2781.500 1958.530 ;
        RECT 14.380 1927.630 2781.500 1939.930 ;
        RECT 14.380 1908.790 2781.500 1921.330 ;
        RECT 14.380 1874.830 2781.500 1902.490 ;
        RECT 14.380 1856.230 2781.500 1868.530 ;
        RECT 14.380 1837.630 2781.500 1849.930 ;
        RECT 14.380 1818.790 2781.500 1831.330 ;
        RECT 14.380 1784.830 2781.500 1812.490 ;
        RECT 14.380 1766.230 2781.500 1778.530 ;
        RECT 14.380 1747.630 2781.500 1759.930 ;
        RECT 14.380 1728.790 2781.500 1741.330 ;
        RECT 14.380 1694.830 2781.500 1722.490 ;
        RECT 14.380 1676.230 2781.500 1688.530 ;
        RECT 14.380 1657.630 2781.500 1669.930 ;
        RECT 14.380 1638.790 2781.500 1651.330 ;
        RECT 14.380 1604.830 2781.500 1632.490 ;
        RECT 14.380 1586.230 2781.500 1598.530 ;
        RECT 14.380 1567.630 2781.500 1579.930 ;
        RECT 14.380 1548.790 2781.500 1561.330 ;
        RECT 14.380 1514.830 2781.500 1542.490 ;
        RECT 14.380 1496.230 2781.500 1508.530 ;
        RECT 14.380 1477.630 2781.500 1489.930 ;
        RECT 14.380 1458.790 2781.500 1471.330 ;
        RECT 14.380 1424.830 2781.500 1452.490 ;
        RECT 14.380 1406.230 2781.500 1418.530 ;
        RECT 14.380 1387.630 2781.500 1399.930 ;
        RECT 14.380 1368.790 2781.500 1381.330 ;
        RECT 14.380 1334.830 2781.500 1362.490 ;
        RECT 14.380 1316.230 2781.500 1328.530 ;
        RECT 14.380 1297.630 2781.500 1309.930 ;
        RECT 14.380 1278.790 2781.500 1291.330 ;
        RECT 14.380 1244.830 2781.500 1272.490 ;
        RECT 14.380 1226.230 2781.500 1238.530 ;
        RECT 14.380 1207.630 2781.500 1219.930 ;
        RECT 14.380 1188.790 2781.500 1201.330 ;
        RECT 14.380 1154.830 2781.500 1182.490 ;
        RECT 14.380 1136.230 2781.500 1148.530 ;
        RECT 14.380 1117.630 2781.500 1129.930 ;
        RECT 14.380 1098.790 2781.500 1111.330 ;
        RECT 14.380 1064.830 2781.500 1092.490 ;
        RECT 14.380 1046.230 2781.500 1058.530 ;
        RECT 14.380 1027.630 2781.500 1039.930 ;
        RECT 14.380 1008.790 2781.500 1021.330 ;
        RECT 14.380 974.830 2781.500 1002.490 ;
        RECT 14.380 956.230 2781.500 968.530 ;
        RECT 14.380 937.630 2781.500 949.930 ;
        RECT 14.380 918.790 2781.500 931.330 ;
        RECT 14.380 884.830 2781.500 912.490 ;
        RECT 14.380 866.230 2781.500 878.530 ;
        RECT 14.380 847.630 2781.500 859.930 ;
        RECT 14.380 828.790 2781.500 841.330 ;
        RECT 14.380 794.830 2781.500 822.490 ;
        RECT 14.380 776.230 2781.500 788.530 ;
        RECT 14.380 757.630 2781.500 769.930 ;
        RECT 14.380 738.790 2781.500 751.330 ;
        RECT 14.380 704.830 2781.500 732.490 ;
        RECT 14.380 686.230 2781.500 698.530 ;
        RECT 14.380 667.630 2781.500 679.930 ;
        RECT 14.380 648.790 2781.500 661.330 ;
        RECT 14.380 614.830 2781.500 642.490 ;
        RECT 14.380 596.230 2781.500 608.530 ;
        RECT 14.380 577.630 2781.500 589.930 ;
        RECT 14.380 558.790 2781.500 571.330 ;
        RECT 14.380 524.830 2781.500 552.490 ;
        RECT 14.380 506.230 2781.500 518.530 ;
        RECT 14.380 487.630 2781.500 499.930 ;
        RECT 14.380 468.790 2781.500 481.330 ;
        RECT 14.380 434.830 2781.500 462.490 ;
        RECT 14.380 416.230 2781.500 428.530 ;
        RECT 14.380 397.630 2781.500 409.930 ;
        RECT 14.380 378.790 2781.500 391.330 ;
        RECT 14.380 344.830 2781.500 372.490 ;
        RECT 14.380 326.230 2781.500 338.530 ;
        RECT 14.380 307.630 2781.500 319.930 ;
        RECT 14.380 288.790 2781.500 301.330 ;
        RECT 14.380 254.830 2781.500 282.490 ;
        RECT 14.380 236.230 2781.500 248.530 ;
        RECT 14.380 217.630 2781.500 229.930 ;
        RECT 14.380 198.790 2781.500 211.330 ;
        RECT 14.380 164.830 2781.500 192.490 ;
        RECT 14.380 146.230 2781.500 158.530 ;
        RECT 14.380 127.630 2781.500 139.930 ;
        RECT 14.380 108.790 2781.500 121.330 ;
        RECT 14.380 74.830 2781.500 102.490 ;
        RECT 14.380 56.230 2781.500 68.530 ;
        RECT 14.380 38.300 2781.500 49.930 ;
  END
END user_project_wrapper
END LIBRARY

