magic
tech sky130A
magscale 1 2
timestamp 1654573858
<< obsli1 >>
rect 552 527 234140 19601
<< obsm1 >>
rect 198 76 234140 36712
<< metal2 >>
rect 846 36688 902 37088
rect 2594 36688 2650 37088
rect 4434 36688 4490 37088
rect 6274 36688 6330 37088
rect 8114 36688 8170 37088
rect 9954 36688 10010 37088
rect 11794 36688 11850 37088
rect 13634 36688 13690 37088
rect 15474 36688 15530 37088
rect 17314 36688 17370 37088
rect 19154 36688 19210 37088
rect 20994 36688 21050 37088
rect 22834 36688 22890 37088
rect 24674 36688 24730 37088
rect 26514 36688 26570 37088
rect 28262 36688 28318 37088
rect 30102 36688 30158 37088
rect 31942 36688 31998 37088
rect 33782 36688 33838 37088
rect 35622 36688 35678 37088
rect 37462 36688 37518 37088
rect 39302 36688 39358 37088
rect 41142 36688 41198 37088
rect 42982 36688 43038 37088
rect 44822 36688 44878 37088
rect 46662 36688 46718 37088
rect 48502 36688 48558 37088
rect 50342 36688 50398 37088
rect 52182 36688 52238 37088
rect 53930 36688 53986 37088
rect 55770 36688 55826 37088
rect 57610 36688 57666 37088
rect 59450 36688 59506 37088
rect 61290 36688 61346 37088
rect 63130 36688 63186 37088
rect 64970 36688 65026 37088
rect 66810 36688 66866 37088
rect 68650 36688 68706 37088
rect 70490 36688 70546 37088
rect 72330 36688 72386 37088
rect 74170 36688 74226 37088
rect 76010 36688 76066 37088
rect 77850 36688 77906 37088
rect 79598 36688 79654 37088
rect 81438 36688 81494 37088
rect 83278 36688 83334 37088
rect 85118 36688 85174 37088
rect 86958 36688 87014 37088
rect 88798 36688 88854 37088
rect 90638 36688 90694 37088
rect 92478 36688 92534 37088
rect 94318 36688 94374 37088
rect 96158 36688 96214 37088
rect 97998 36688 98054 37088
rect 99838 36688 99894 37088
rect 101678 36688 101734 37088
rect 103518 36688 103574 37088
rect 105266 36688 105322 37088
rect 107106 36688 107162 37088
rect 108946 36688 109002 37088
rect 110786 36688 110842 37088
rect 112626 36688 112682 37088
rect 114466 36688 114522 37088
rect 116306 36688 116362 37088
rect 118146 36688 118202 37088
rect 119986 36688 120042 37088
rect 121826 36688 121882 37088
rect 123666 36688 123722 37088
rect 125506 36688 125562 37088
rect 127346 36688 127402 37088
rect 129186 36688 129242 37088
rect 131026 36688 131082 37088
rect 132774 36688 132830 37088
rect 134614 36688 134670 37088
rect 136454 36688 136510 37088
rect 138294 36688 138350 37088
rect 140134 36688 140190 37088
rect 141974 36688 142030 37088
rect 143814 36688 143870 37088
rect 145654 36688 145710 37088
rect 147494 36688 147550 37088
rect 149334 36688 149390 37088
rect 151174 36688 151230 37088
rect 153014 36688 153070 37088
rect 154854 36688 154910 37088
rect 156694 36688 156750 37088
rect 158442 36688 158498 37088
rect 160282 36688 160338 37088
rect 162122 36688 162178 37088
rect 163962 36688 164018 37088
rect 165802 36688 165858 37088
rect 167642 36688 167698 37088
rect 169482 36688 169538 37088
rect 171322 36688 171378 37088
rect 173162 36688 173218 37088
rect 175002 36688 175058 37088
rect 176842 36688 176898 37088
rect 178682 36688 178738 37088
rect 180522 36688 180578 37088
rect 182362 36688 182418 37088
rect 184110 36688 184166 37088
rect 185950 36688 186006 37088
rect 187790 36688 187846 37088
rect 189630 36688 189686 37088
rect 191470 36688 191526 37088
rect 193310 36688 193366 37088
rect 195150 36688 195206 37088
rect 196990 36688 197046 37088
rect 198830 36688 198886 37088
rect 200670 36688 200726 37088
rect 202510 36688 202566 37088
rect 204350 36688 204406 37088
rect 206190 36688 206246 37088
rect 208030 36688 208086 37088
rect 209778 36688 209834 37088
rect 211618 36688 211674 37088
rect 213458 36688 213514 37088
rect 215298 36688 215354 37088
rect 217138 36688 217194 37088
rect 218978 36688 219034 37088
rect 220818 36688 220874 37088
rect 222658 36688 222714 37088
rect 224498 36688 224554 37088
rect 226338 36688 226394 37088
rect 228178 36688 228234 37088
rect 230018 36688 230074 37088
rect 231858 36688 231914 37088
rect 233698 36688 233754 37088
rect 1766 0 1822 400
rect 5354 0 5410 400
rect 9034 0 9090 400
rect 12714 0 12770 400
rect 16394 0 16450 400
rect 20074 0 20130 400
rect 23754 0 23810 400
rect 27434 0 27490 400
rect 31022 0 31078 400
rect 34702 0 34758 400
rect 38382 0 38438 400
rect 42062 0 42118 400
rect 45742 0 45798 400
rect 49422 0 49478 400
rect 53102 0 53158 400
rect 56690 0 56746 400
rect 60370 0 60426 400
rect 64050 0 64106 400
rect 67730 0 67786 400
rect 71410 0 71466 400
rect 75090 0 75146 400
rect 78770 0 78826 400
rect 82358 0 82414 400
rect 86038 0 86094 400
rect 89718 0 89774 400
rect 93398 0 93454 400
rect 97078 0 97134 400
rect 100758 0 100814 400
rect 104438 0 104494 400
rect 108026 0 108082 400
rect 111706 0 111762 400
rect 115386 0 115442 400
rect 119066 0 119122 400
rect 122746 0 122802 400
rect 126426 0 126482 400
rect 130106 0 130162 400
rect 133694 0 133750 400
rect 137374 0 137430 400
rect 141054 0 141110 400
rect 144734 0 144790 400
rect 148414 0 148470 400
rect 152094 0 152150 400
rect 155774 0 155830 400
rect 159362 0 159418 400
rect 163042 0 163098 400
rect 166722 0 166778 400
rect 170402 0 170458 400
rect 174082 0 174138 400
rect 177762 0 177818 400
rect 181442 0 181498 400
rect 185030 0 185086 400
rect 188710 0 188766 400
rect 192390 0 192446 400
rect 196070 0 196126 400
rect 199750 0 199806 400
rect 203430 0 203486 400
rect 207110 0 207166 400
rect 210698 0 210754 400
rect 214378 0 214434 400
rect 218058 0 218114 400
rect 221738 0 221794 400
rect 225418 0 225474 400
rect 229098 0 229154 400
rect 232778 0 232834 400
<< obsm2 >>
rect 204 36632 790 36802
rect 958 36632 2538 36802
rect 2706 36632 4378 36802
rect 4546 36632 6218 36802
rect 6386 36632 8058 36802
rect 8226 36632 9898 36802
rect 10066 36632 11738 36802
rect 11906 36632 13578 36802
rect 13746 36632 15418 36802
rect 15586 36632 17258 36802
rect 17426 36632 19098 36802
rect 19266 36632 20938 36802
rect 21106 36632 22778 36802
rect 22946 36632 24618 36802
rect 24786 36632 26458 36802
rect 26626 36632 28206 36802
rect 28374 36632 30046 36802
rect 30214 36632 31886 36802
rect 32054 36632 33726 36802
rect 33894 36632 35566 36802
rect 35734 36632 37406 36802
rect 37574 36632 39246 36802
rect 39414 36632 41086 36802
rect 41254 36632 42926 36802
rect 43094 36632 44766 36802
rect 44934 36632 46606 36802
rect 46774 36632 48446 36802
rect 48614 36632 50286 36802
rect 50454 36632 52126 36802
rect 52294 36632 53874 36802
rect 54042 36632 55714 36802
rect 55882 36632 57554 36802
rect 57722 36632 59394 36802
rect 59562 36632 61234 36802
rect 61402 36632 63074 36802
rect 63242 36632 64914 36802
rect 65082 36632 66754 36802
rect 66922 36632 68594 36802
rect 68762 36632 70434 36802
rect 70602 36632 72274 36802
rect 72442 36632 74114 36802
rect 74282 36632 75954 36802
rect 76122 36632 77794 36802
rect 77962 36632 79542 36802
rect 79710 36632 81382 36802
rect 81550 36632 83222 36802
rect 83390 36632 85062 36802
rect 85230 36632 86902 36802
rect 87070 36632 88742 36802
rect 88910 36632 90582 36802
rect 90750 36632 92422 36802
rect 92590 36632 94262 36802
rect 94430 36632 96102 36802
rect 96270 36632 97942 36802
rect 98110 36632 99782 36802
rect 99950 36632 101622 36802
rect 101790 36632 103462 36802
rect 103630 36632 105210 36802
rect 105378 36632 107050 36802
rect 107218 36632 108890 36802
rect 109058 36632 110730 36802
rect 110898 36632 112570 36802
rect 112738 36632 114410 36802
rect 114578 36632 116250 36802
rect 116418 36632 118090 36802
rect 118258 36632 119930 36802
rect 120098 36632 121770 36802
rect 121938 36632 123610 36802
rect 123778 36632 125450 36802
rect 125618 36632 127290 36802
rect 127458 36632 129130 36802
rect 129298 36632 130970 36802
rect 131138 36632 132718 36802
rect 132886 36632 134558 36802
rect 134726 36632 136398 36802
rect 136566 36632 138238 36802
rect 138406 36632 140078 36802
rect 140246 36632 141918 36802
rect 142086 36632 143758 36802
rect 143926 36632 145598 36802
rect 145766 36632 147438 36802
rect 147606 36632 149278 36802
rect 149446 36632 151118 36802
rect 151286 36632 152958 36802
rect 153126 36632 154798 36802
rect 154966 36632 156638 36802
rect 156806 36632 158386 36802
rect 158554 36632 160226 36802
rect 160394 36632 162066 36802
rect 162234 36632 163906 36802
rect 164074 36632 165746 36802
rect 165914 36632 167586 36802
rect 167754 36632 169426 36802
rect 169594 36632 171266 36802
rect 171434 36632 173106 36802
rect 173274 36632 174946 36802
rect 175114 36632 176786 36802
rect 176954 36632 178626 36802
rect 178794 36632 180466 36802
rect 180634 36632 182306 36802
rect 182474 36632 184054 36802
rect 184222 36632 185894 36802
rect 186062 36632 187734 36802
rect 187902 36632 189574 36802
rect 189742 36632 191414 36802
rect 191582 36632 193254 36802
rect 193422 36632 195094 36802
rect 195262 36632 196934 36802
rect 197102 36632 198774 36802
rect 198942 36632 200614 36802
rect 200782 36632 202454 36802
rect 202622 36632 204294 36802
rect 204462 36632 206134 36802
rect 206302 36632 207974 36802
rect 208142 36632 209722 36802
rect 209890 36632 211562 36802
rect 211730 36632 213402 36802
rect 213570 36632 215242 36802
rect 215410 36632 217082 36802
rect 217250 36632 218922 36802
rect 219090 36632 220762 36802
rect 220930 36632 222602 36802
rect 222770 36632 224442 36802
rect 224610 36632 226282 36802
rect 226450 36632 228122 36802
rect 228290 36632 229962 36802
rect 230130 36632 231802 36802
rect 231970 36632 233642 36802
rect 233810 36632 233936 36802
rect 204 456 233936 36632
rect 204 31 1710 456
rect 1878 31 5298 456
rect 5466 31 8978 456
rect 9146 31 12658 456
rect 12826 31 16338 456
rect 16506 31 20018 456
rect 20186 31 23698 456
rect 23866 31 27378 456
rect 27546 31 30966 456
rect 31134 31 34646 456
rect 34814 31 38326 456
rect 38494 31 42006 456
rect 42174 31 45686 456
rect 45854 31 49366 456
rect 49534 31 53046 456
rect 53214 31 56634 456
rect 56802 31 60314 456
rect 60482 31 63994 456
rect 64162 31 67674 456
rect 67842 31 71354 456
rect 71522 31 75034 456
rect 75202 31 78714 456
rect 78882 31 82302 456
rect 82470 31 85982 456
rect 86150 31 89662 456
rect 89830 31 93342 456
rect 93510 31 97022 456
rect 97190 31 100702 456
rect 100870 31 104382 456
rect 104550 31 107970 456
rect 108138 31 111650 456
rect 111818 31 115330 456
rect 115498 31 119010 456
rect 119178 31 122690 456
rect 122858 31 126370 456
rect 126538 31 130050 456
rect 130218 31 133638 456
rect 133806 31 137318 456
rect 137486 31 140998 456
rect 141166 31 144678 456
rect 144846 31 148358 456
rect 148526 31 152038 456
rect 152206 31 155718 456
rect 155886 31 159306 456
rect 159474 31 162986 456
rect 163154 31 166666 456
rect 166834 31 170346 456
rect 170514 31 174026 456
rect 174194 31 177706 456
rect 177874 31 181386 456
rect 181554 31 184974 456
rect 185142 31 188654 456
rect 188822 31 192334 456
rect 192502 31 196014 456
rect 196182 31 199694 456
rect 199862 31 203374 456
rect 203542 31 207054 456
rect 207222 31 210642 456
rect 210810 31 214322 456
rect 214490 31 218002 456
rect 218170 31 221682 456
rect 221850 31 225362 456
rect 225530 31 229042 456
rect 229210 31 232722 456
rect 232890 31 233936 456
<< metal3 >>
rect 234292 35640 234692 35760
rect 0 34416 400 34536
rect 234292 33056 234692 33176
rect 234292 30336 234692 30456
rect 0 29112 400 29232
rect 234292 27752 234692 27872
rect 234292 25032 234692 25152
rect 0 23808 400 23928
rect 234292 22448 234692 22568
rect 234292 19728 234692 19848
rect 0 18504 400 18624
rect 234292 17144 234692 17264
rect 234292 14424 234692 14544
rect 0 13200 400 13320
rect 234292 11840 234692 11960
rect 234292 9120 234692 9240
rect 0 7896 400 8016
rect 234292 6536 234692 6656
rect 234292 3816 234692 3936
rect 0 2592 400 2712
rect 234292 1232 234692 1352
<< obsm3 >>
rect 381 35840 234292 36481
rect 381 35560 234212 35840
rect 381 34616 234292 35560
rect 480 34336 234292 34616
rect 381 33256 234292 34336
rect 381 32976 234212 33256
rect 381 30536 234292 32976
rect 381 30256 234212 30536
rect 381 29312 234292 30256
rect 480 29032 234292 29312
rect 381 27952 234292 29032
rect 381 27672 234212 27952
rect 381 25232 234292 27672
rect 381 24952 234212 25232
rect 381 24008 234292 24952
rect 480 23728 234292 24008
rect 381 22648 234292 23728
rect 381 22368 234212 22648
rect 381 19928 234292 22368
rect 381 19648 234212 19928
rect 381 18704 234292 19648
rect 480 18424 234292 18704
rect 381 17344 234292 18424
rect 381 17064 234212 17344
rect 381 14624 234292 17064
rect 381 14344 234212 14624
rect 381 13400 234292 14344
rect 480 13120 234292 13400
rect 381 12040 234292 13120
rect 381 11760 234212 12040
rect 381 9320 234292 11760
rect 381 9040 234212 9320
rect 381 8096 234292 9040
rect 480 7816 234292 8096
rect 381 6736 234292 7816
rect 381 6456 234212 6736
rect 381 4016 234292 6456
rect 381 3736 234212 4016
rect 381 2792 234292 3736
rect 480 2512 234292 2792
rect 381 1432 234292 2512
rect 381 1152 234212 1432
rect 381 35 234292 1152
<< metal4 >>
rect 1242 496 1862 36496
rect 19242 496 19862 36496
rect 37242 496 37862 36496
rect 55242 496 55862 36496
rect 73242 496 73862 36496
rect 91242 496 91862 36496
rect 109242 496 109862 36496
rect 127242 496 127862 36496
rect 145242 496 145862 36496
rect 163242 496 163862 36496
rect 181242 496 181862 36496
rect 199242 496 199862 36496
rect 217242 496 217862 36496
<< obsm4 >>
rect 979 416 1162 35597
rect 1942 416 19162 35597
rect 19942 416 37162 35597
rect 37942 416 55162 35597
rect 55942 416 73162 35597
rect 73942 416 91162 35597
rect 91942 416 109162 35597
rect 109942 416 127162 35597
rect 127942 416 145162 35597
rect 145942 416 163162 35597
rect 163942 416 181162 35597
rect 181942 416 199162 35597
rect 199942 416 215589 35597
rect 979 171 215589 416
<< labels >>
rlabel metal3 s 234292 25032 234692 25152 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 234292 27752 234692 27872 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 234292 30336 234692 30456 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 234292 33056 234692 33176 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 234292 35640 234692 35760 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 0 7896 400 8016 6 A1[0]
port 6 nsew signal input
rlabel metal3 s 0 13200 400 13320 6 A1[1]
port 7 nsew signal input
rlabel metal3 s 0 18504 400 18624 6 A1[2]
port 8 nsew signal input
rlabel metal3 s 0 23808 400 23928 6 A1[3]
port 9 nsew signal input
rlabel metal3 s 0 29112 400 29232 6 A1[4]
port 10 nsew signal input
rlabel metal3 s 0 2592 400 2712 6 CLK
port 11 nsew signal input
rlabel metal2 s 1766 0 1822 400 6 Di0[0]
port 12 nsew signal input
rlabel metal2 s 38382 0 38438 400 6 Di0[10]
port 13 nsew signal input
rlabel metal2 s 42062 0 42118 400 6 Di0[11]
port 14 nsew signal input
rlabel metal2 s 45742 0 45798 400 6 Di0[12]
port 15 nsew signal input
rlabel metal2 s 49422 0 49478 400 6 Di0[13]
port 16 nsew signal input
rlabel metal2 s 53102 0 53158 400 6 Di0[14]
port 17 nsew signal input
rlabel metal2 s 56690 0 56746 400 6 Di0[15]
port 18 nsew signal input
rlabel metal2 s 60370 0 60426 400 6 Di0[16]
port 19 nsew signal input
rlabel metal2 s 64050 0 64106 400 6 Di0[17]
port 20 nsew signal input
rlabel metal2 s 67730 0 67786 400 6 Di0[18]
port 21 nsew signal input
rlabel metal2 s 71410 0 71466 400 6 Di0[19]
port 22 nsew signal input
rlabel metal2 s 5354 0 5410 400 6 Di0[1]
port 23 nsew signal input
rlabel metal2 s 75090 0 75146 400 6 Di0[20]
port 24 nsew signal input
rlabel metal2 s 78770 0 78826 400 6 Di0[21]
port 25 nsew signal input
rlabel metal2 s 82358 0 82414 400 6 Di0[22]
port 26 nsew signal input
rlabel metal2 s 86038 0 86094 400 6 Di0[23]
port 27 nsew signal input
rlabel metal2 s 89718 0 89774 400 6 Di0[24]
port 28 nsew signal input
rlabel metal2 s 93398 0 93454 400 6 Di0[25]
port 29 nsew signal input
rlabel metal2 s 97078 0 97134 400 6 Di0[26]
port 30 nsew signal input
rlabel metal2 s 100758 0 100814 400 6 Di0[27]
port 31 nsew signal input
rlabel metal2 s 104438 0 104494 400 6 Di0[28]
port 32 nsew signal input
rlabel metal2 s 108026 0 108082 400 6 Di0[29]
port 33 nsew signal input
rlabel metal2 s 9034 0 9090 400 6 Di0[2]
port 34 nsew signal input
rlabel metal2 s 111706 0 111762 400 6 Di0[30]
port 35 nsew signal input
rlabel metal2 s 115386 0 115442 400 6 Di0[31]
port 36 nsew signal input
rlabel metal2 s 119066 0 119122 400 6 Di0[32]
port 37 nsew signal input
rlabel metal2 s 122746 0 122802 400 6 Di0[33]
port 38 nsew signal input
rlabel metal2 s 126426 0 126482 400 6 Di0[34]
port 39 nsew signal input
rlabel metal2 s 130106 0 130162 400 6 Di0[35]
port 40 nsew signal input
rlabel metal2 s 133694 0 133750 400 6 Di0[36]
port 41 nsew signal input
rlabel metal2 s 137374 0 137430 400 6 Di0[37]
port 42 nsew signal input
rlabel metal2 s 141054 0 141110 400 6 Di0[38]
port 43 nsew signal input
rlabel metal2 s 144734 0 144790 400 6 Di0[39]
port 44 nsew signal input
rlabel metal2 s 12714 0 12770 400 6 Di0[3]
port 45 nsew signal input
rlabel metal2 s 148414 0 148470 400 6 Di0[40]
port 46 nsew signal input
rlabel metal2 s 152094 0 152150 400 6 Di0[41]
port 47 nsew signal input
rlabel metal2 s 155774 0 155830 400 6 Di0[42]
port 48 nsew signal input
rlabel metal2 s 159362 0 159418 400 6 Di0[43]
port 49 nsew signal input
rlabel metal2 s 163042 0 163098 400 6 Di0[44]
port 50 nsew signal input
rlabel metal2 s 166722 0 166778 400 6 Di0[45]
port 51 nsew signal input
rlabel metal2 s 170402 0 170458 400 6 Di0[46]
port 52 nsew signal input
rlabel metal2 s 174082 0 174138 400 6 Di0[47]
port 53 nsew signal input
rlabel metal2 s 177762 0 177818 400 6 Di0[48]
port 54 nsew signal input
rlabel metal2 s 181442 0 181498 400 6 Di0[49]
port 55 nsew signal input
rlabel metal2 s 16394 0 16450 400 6 Di0[4]
port 56 nsew signal input
rlabel metal2 s 185030 0 185086 400 6 Di0[50]
port 57 nsew signal input
rlabel metal2 s 188710 0 188766 400 6 Di0[51]
port 58 nsew signal input
rlabel metal2 s 192390 0 192446 400 6 Di0[52]
port 59 nsew signal input
rlabel metal2 s 196070 0 196126 400 6 Di0[53]
port 60 nsew signal input
rlabel metal2 s 199750 0 199806 400 6 Di0[54]
port 61 nsew signal input
rlabel metal2 s 203430 0 203486 400 6 Di0[55]
port 62 nsew signal input
rlabel metal2 s 207110 0 207166 400 6 Di0[56]
port 63 nsew signal input
rlabel metal2 s 210698 0 210754 400 6 Di0[57]
port 64 nsew signal input
rlabel metal2 s 214378 0 214434 400 6 Di0[58]
port 65 nsew signal input
rlabel metal2 s 218058 0 218114 400 6 Di0[59]
port 66 nsew signal input
rlabel metal2 s 20074 0 20130 400 6 Di0[5]
port 67 nsew signal input
rlabel metal2 s 221738 0 221794 400 6 Di0[60]
port 68 nsew signal input
rlabel metal2 s 225418 0 225474 400 6 Di0[61]
port 69 nsew signal input
rlabel metal2 s 229098 0 229154 400 6 Di0[62]
port 70 nsew signal input
rlabel metal2 s 232778 0 232834 400 6 Di0[63]
port 71 nsew signal input
rlabel metal2 s 23754 0 23810 400 6 Di0[6]
port 72 nsew signal input
rlabel metal2 s 27434 0 27490 400 6 Di0[7]
port 73 nsew signal input
rlabel metal2 s 31022 0 31078 400 6 Di0[8]
port 74 nsew signal input
rlabel metal2 s 34702 0 34758 400 6 Di0[9]
port 75 nsew signal input
rlabel metal2 s 846 36688 902 37088 6 Do0[0]
port 76 nsew signal output
rlabel metal2 s 19154 36688 19210 37088 6 Do0[10]
port 77 nsew signal output
rlabel metal2 s 22834 36688 22890 37088 6 Do0[11]
port 78 nsew signal output
rlabel metal2 s 26514 36688 26570 37088 6 Do0[12]
port 79 nsew signal output
rlabel metal2 s 30102 36688 30158 37088 6 Do0[13]
port 80 nsew signal output
rlabel metal2 s 33782 36688 33838 37088 6 Do0[14]
port 81 nsew signal output
rlabel metal2 s 37462 36688 37518 37088 6 Do0[15]
port 82 nsew signal output
rlabel metal2 s 41142 36688 41198 37088 6 Do0[16]
port 83 nsew signal output
rlabel metal2 s 44822 36688 44878 37088 6 Do0[17]
port 84 nsew signal output
rlabel metal2 s 48502 36688 48558 37088 6 Do0[18]
port 85 nsew signal output
rlabel metal2 s 52182 36688 52238 37088 6 Do0[19]
port 86 nsew signal output
rlabel metal2 s 2594 36688 2650 37088 6 Do0[1]
port 87 nsew signal output
rlabel metal2 s 55770 36688 55826 37088 6 Do0[20]
port 88 nsew signal output
rlabel metal2 s 57610 36688 57666 37088 6 Do0[21]
port 89 nsew signal output
rlabel metal2 s 59450 36688 59506 37088 6 Do0[22]
port 90 nsew signal output
rlabel metal2 s 61290 36688 61346 37088 6 Do0[23]
port 91 nsew signal output
rlabel metal2 s 63130 36688 63186 37088 6 Do0[24]
port 92 nsew signal output
rlabel metal2 s 64970 36688 65026 37088 6 Do0[25]
port 93 nsew signal output
rlabel metal2 s 66810 36688 66866 37088 6 Do0[26]
port 94 nsew signal output
rlabel metal2 s 68650 36688 68706 37088 6 Do0[27]
port 95 nsew signal output
rlabel metal2 s 70490 36688 70546 37088 6 Do0[28]
port 96 nsew signal output
rlabel metal2 s 72330 36688 72386 37088 6 Do0[29]
port 97 nsew signal output
rlabel metal2 s 4434 36688 4490 37088 6 Do0[2]
port 98 nsew signal output
rlabel metal2 s 74170 36688 74226 37088 6 Do0[30]
port 99 nsew signal output
rlabel metal2 s 76010 36688 76066 37088 6 Do0[31]
port 100 nsew signal output
rlabel metal2 s 77850 36688 77906 37088 6 Do0[32]
port 101 nsew signal output
rlabel metal2 s 79598 36688 79654 37088 6 Do0[33]
port 102 nsew signal output
rlabel metal2 s 81438 36688 81494 37088 6 Do0[34]
port 103 nsew signal output
rlabel metal2 s 83278 36688 83334 37088 6 Do0[35]
port 104 nsew signal output
rlabel metal2 s 85118 36688 85174 37088 6 Do0[36]
port 105 nsew signal output
rlabel metal2 s 86958 36688 87014 37088 6 Do0[37]
port 106 nsew signal output
rlabel metal2 s 88798 36688 88854 37088 6 Do0[38]
port 107 nsew signal output
rlabel metal2 s 90638 36688 90694 37088 6 Do0[39]
port 108 nsew signal output
rlabel metal2 s 6274 36688 6330 37088 6 Do0[3]
port 109 nsew signal output
rlabel metal2 s 92478 36688 92534 37088 6 Do0[40]
port 110 nsew signal output
rlabel metal2 s 94318 36688 94374 37088 6 Do0[41]
port 111 nsew signal output
rlabel metal2 s 96158 36688 96214 37088 6 Do0[42]
port 112 nsew signal output
rlabel metal2 s 97998 36688 98054 37088 6 Do0[43]
port 113 nsew signal output
rlabel metal2 s 99838 36688 99894 37088 6 Do0[44]
port 114 nsew signal output
rlabel metal2 s 101678 36688 101734 37088 6 Do0[45]
port 115 nsew signal output
rlabel metal2 s 103518 36688 103574 37088 6 Do0[46]
port 116 nsew signal output
rlabel metal2 s 105266 36688 105322 37088 6 Do0[47]
port 117 nsew signal output
rlabel metal2 s 107106 36688 107162 37088 6 Do0[48]
port 118 nsew signal output
rlabel metal2 s 108946 36688 109002 37088 6 Do0[49]
port 119 nsew signal output
rlabel metal2 s 8114 36688 8170 37088 6 Do0[4]
port 120 nsew signal output
rlabel metal2 s 110786 36688 110842 37088 6 Do0[50]
port 121 nsew signal output
rlabel metal2 s 112626 36688 112682 37088 6 Do0[51]
port 122 nsew signal output
rlabel metal2 s 114466 36688 114522 37088 6 Do0[52]
port 123 nsew signal output
rlabel metal2 s 116306 36688 116362 37088 6 Do0[53]
port 124 nsew signal output
rlabel metal2 s 118146 36688 118202 37088 6 Do0[54]
port 125 nsew signal output
rlabel metal2 s 119986 36688 120042 37088 6 Do0[55]
port 126 nsew signal output
rlabel metal2 s 121826 36688 121882 37088 6 Do0[56]
port 127 nsew signal output
rlabel metal2 s 123666 36688 123722 37088 6 Do0[57]
port 128 nsew signal output
rlabel metal2 s 125506 36688 125562 37088 6 Do0[58]
port 129 nsew signal output
rlabel metal2 s 127346 36688 127402 37088 6 Do0[59]
port 130 nsew signal output
rlabel metal2 s 9954 36688 10010 37088 6 Do0[5]
port 131 nsew signal output
rlabel metal2 s 129186 36688 129242 37088 6 Do0[60]
port 132 nsew signal output
rlabel metal2 s 131026 36688 131082 37088 6 Do0[61]
port 133 nsew signal output
rlabel metal2 s 132774 36688 132830 37088 6 Do0[62]
port 134 nsew signal output
rlabel metal2 s 134614 36688 134670 37088 6 Do0[63]
port 135 nsew signal output
rlabel metal2 s 11794 36688 11850 37088 6 Do0[6]
port 136 nsew signal output
rlabel metal2 s 13634 36688 13690 37088 6 Do0[7]
port 137 nsew signal output
rlabel metal2 s 15474 36688 15530 37088 6 Do0[8]
port 138 nsew signal output
rlabel metal2 s 17314 36688 17370 37088 6 Do0[9]
port 139 nsew signal output
rlabel metal2 s 20994 36688 21050 37088 6 Do1[0]
port 140 nsew signal output
rlabel metal2 s 136454 36688 136510 37088 6 Do1[10]
port 141 nsew signal output
rlabel metal2 s 138294 36688 138350 37088 6 Do1[11]
port 142 nsew signal output
rlabel metal2 s 140134 36688 140190 37088 6 Do1[12]
port 143 nsew signal output
rlabel metal2 s 141974 36688 142030 37088 6 Do1[13]
port 144 nsew signal output
rlabel metal2 s 143814 36688 143870 37088 6 Do1[14]
port 145 nsew signal output
rlabel metal2 s 145654 36688 145710 37088 6 Do1[15]
port 146 nsew signal output
rlabel metal2 s 147494 36688 147550 37088 6 Do1[16]
port 147 nsew signal output
rlabel metal2 s 149334 36688 149390 37088 6 Do1[17]
port 148 nsew signal output
rlabel metal2 s 151174 36688 151230 37088 6 Do1[18]
port 149 nsew signal output
rlabel metal2 s 153014 36688 153070 37088 6 Do1[19]
port 150 nsew signal output
rlabel metal2 s 24674 36688 24730 37088 6 Do1[1]
port 151 nsew signal output
rlabel metal2 s 154854 36688 154910 37088 6 Do1[20]
port 152 nsew signal output
rlabel metal2 s 156694 36688 156750 37088 6 Do1[21]
port 153 nsew signal output
rlabel metal2 s 158442 36688 158498 37088 6 Do1[22]
port 154 nsew signal output
rlabel metal2 s 160282 36688 160338 37088 6 Do1[23]
port 155 nsew signal output
rlabel metal2 s 162122 36688 162178 37088 6 Do1[24]
port 156 nsew signal output
rlabel metal2 s 163962 36688 164018 37088 6 Do1[25]
port 157 nsew signal output
rlabel metal2 s 165802 36688 165858 37088 6 Do1[26]
port 158 nsew signal output
rlabel metal2 s 167642 36688 167698 37088 6 Do1[27]
port 159 nsew signal output
rlabel metal2 s 169482 36688 169538 37088 6 Do1[28]
port 160 nsew signal output
rlabel metal2 s 171322 36688 171378 37088 6 Do1[29]
port 161 nsew signal output
rlabel metal2 s 28262 36688 28318 37088 6 Do1[2]
port 162 nsew signal output
rlabel metal2 s 173162 36688 173218 37088 6 Do1[30]
port 163 nsew signal output
rlabel metal2 s 175002 36688 175058 37088 6 Do1[31]
port 164 nsew signal output
rlabel metal2 s 176842 36688 176898 37088 6 Do1[32]
port 165 nsew signal output
rlabel metal2 s 178682 36688 178738 37088 6 Do1[33]
port 166 nsew signal output
rlabel metal2 s 180522 36688 180578 37088 6 Do1[34]
port 167 nsew signal output
rlabel metal2 s 182362 36688 182418 37088 6 Do1[35]
port 168 nsew signal output
rlabel metal2 s 184110 36688 184166 37088 6 Do1[36]
port 169 nsew signal output
rlabel metal2 s 185950 36688 186006 37088 6 Do1[37]
port 170 nsew signal output
rlabel metal2 s 187790 36688 187846 37088 6 Do1[38]
port 171 nsew signal output
rlabel metal2 s 189630 36688 189686 37088 6 Do1[39]
port 172 nsew signal output
rlabel metal2 s 31942 36688 31998 37088 6 Do1[3]
port 173 nsew signal output
rlabel metal2 s 191470 36688 191526 37088 6 Do1[40]
port 174 nsew signal output
rlabel metal2 s 193310 36688 193366 37088 6 Do1[41]
port 175 nsew signal output
rlabel metal2 s 195150 36688 195206 37088 6 Do1[42]
port 176 nsew signal output
rlabel metal2 s 196990 36688 197046 37088 6 Do1[43]
port 177 nsew signal output
rlabel metal2 s 198830 36688 198886 37088 6 Do1[44]
port 178 nsew signal output
rlabel metal2 s 200670 36688 200726 37088 6 Do1[45]
port 179 nsew signal output
rlabel metal2 s 202510 36688 202566 37088 6 Do1[46]
port 180 nsew signal output
rlabel metal2 s 204350 36688 204406 37088 6 Do1[47]
port 181 nsew signal output
rlabel metal2 s 206190 36688 206246 37088 6 Do1[48]
port 182 nsew signal output
rlabel metal2 s 208030 36688 208086 37088 6 Do1[49]
port 183 nsew signal output
rlabel metal2 s 35622 36688 35678 37088 6 Do1[4]
port 184 nsew signal output
rlabel metal2 s 209778 36688 209834 37088 6 Do1[50]
port 185 nsew signal output
rlabel metal2 s 211618 36688 211674 37088 6 Do1[51]
port 186 nsew signal output
rlabel metal2 s 213458 36688 213514 37088 6 Do1[52]
port 187 nsew signal output
rlabel metal2 s 215298 36688 215354 37088 6 Do1[53]
port 188 nsew signal output
rlabel metal2 s 217138 36688 217194 37088 6 Do1[54]
port 189 nsew signal output
rlabel metal2 s 218978 36688 219034 37088 6 Do1[55]
port 190 nsew signal output
rlabel metal2 s 220818 36688 220874 37088 6 Do1[56]
port 191 nsew signal output
rlabel metal2 s 222658 36688 222714 37088 6 Do1[57]
port 192 nsew signal output
rlabel metal2 s 224498 36688 224554 37088 6 Do1[58]
port 193 nsew signal output
rlabel metal2 s 226338 36688 226394 37088 6 Do1[59]
port 194 nsew signal output
rlabel metal2 s 39302 36688 39358 37088 6 Do1[5]
port 195 nsew signal output
rlabel metal2 s 228178 36688 228234 37088 6 Do1[60]
port 196 nsew signal output
rlabel metal2 s 230018 36688 230074 37088 6 Do1[61]
port 197 nsew signal output
rlabel metal2 s 231858 36688 231914 37088 6 Do1[62]
port 198 nsew signal output
rlabel metal2 s 233698 36688 233754 37088 6 Do1[63]
port 199 nsew signal output
rlabel metal2 s 42982 36688 43038 37088 6 Do1[6]
port 200 nsew signal output
rlabel metal2 s 46662 36688 46718 37088 6 Do1[7]
port 201 nsew signal output
rlabel metal2 s 50342 36688 50398 37088 6 Do1[8]
port 202 nsew signal output
rlabel metal2 s 53930 36688 53986 37088 6 Do1[9]
port 203 nsew signal output
rlabel metal3 s 234292 1232 234692 1352 6 EN0
port 204 nsew signal input
rlabel metal3 s 0 34416 400 34536 6 EN1
port 205 nsew signal input
rlabel metal4 s 19242 496 19862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 55242 496 55862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 91242 496 91862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 127242 496 127862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 163242 496 163862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 199242 496 199862 36496 6 VGND
port 206 nsew ground bidirectional
rlabel metal4 s 1242 496 1862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 37242 496 37862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 73242 496 73862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 109242 496 109862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 145242 496 145862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 181242 496 181862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal4 s 217242 496 217862 36496 6 VPWR
port 207 nsew power bidirectional
rlabel metal3 s 234292 3816 234692 3936 6 WE0[0]
port 208 nsew signal input
rlabel metal3 s 234292 6536 234692 6656 6 WE0[1]
port 209 nsew signal input
rlabel metal3 s 234292 9120 234692 9240 6 WE0[2]
port 210 nsew signal input
rlabel metal3 s 234292 11840 234692 11960 6 WE0[3]
port 211 nsew signal input
rlabel metal3 s 234292 14424 234692 14544 6 WE0[4]
port 212 nsew signal input
rlabel metal3 s 234292 17144 234692 17264 6 WE0[5]
port 213 nsew signal input
rlabel metal3 s 234292 19728 234692 19848 6 WE0[6]
port 214 nsew signal input
rlabel metal3 s 234292 22448 234692 22568 6 WE0[7]
port 215 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 234692 37088
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17778744
string GDS_FILE /mnt/dffram/build/32x64_1RW1R/openlane/runs/RUN_2022.06.07_03.39.53/results/signoff/RAM32_1RW1R.magic.gds
string GDS_START 150134
<< end >>

