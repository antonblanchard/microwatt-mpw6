magic
tech sky130A
magscale 1 2
timestamp 1654578501
<< obsli1 >>
rect 4048 20111 312708 177361
<< obsm1 >>
rect 290 76 316190 197464
<< metal2 >>
rect 2410 197072 2466 197472
rect 7286 197072 7342 197472
rect 12254 197072 12310 197472
rect 17222 197072 17278 197472
rect 22190 197072 22246 197472
rect 27066 197072 27122 197472
rect 32034 197072 32090 197472
rect 37002 197072 37058 197472
rect 41970 197072 42026 197472
rect 46938 197072 46994 197472
rect 51814 197072 51870 197472
rect 56782 197072 56838 197472
rect 61750 197072 61806 197472
rect 66718 197072 66774 197472
rect 71686 197072 71742 197472
rect 76562 197072 76618 197472
rect 81530 197072 81586 197472
rect 86498 197072 86554 197472
rect 91466 197072 91522 197472
rect 96434 197072 96490 197472
rect 101310 197072 101366 197472
rect 106278 197072 106334 197472
rect 111246 197072 111302 197472
rect 116214 197072 116270 197472
rect 121182 197072 121238 197472
rect 126058 197072 126114 197472
rect 131026 197072 131082 197472
rect 135994 197072 136050 197472
rect 140962 197072 141018 197472
rect 145930 197072 145986 197472
rect 150806 197072 150862 197472
rect 155774 197072 155830 197472
rect 160742 197072 160798 197472
rect 165710 197072 165766 197472
rect 170678 197072 170734 197472
rect 175554 197072 175610 197472
rect 180522 197072 180578 197472
rect 185490 197072 185546 197472
rect 190458 197072 190514 197472
rect 195426 197072 195482 197472
rect 200302 197072 200358 197472
rect 205270 197072 205326 197472
rect 210238 197072 210294 197472
rect 215206 197072 215262 197472
rect 220174 197072 220230 197472
rect 225050 197072 225106 197472
rect 230018 197072 230074 197472
rect 234986 197072 235042 197472
rect 239954 197072 240010 197472
rect 244922 197072 244978 197472
rect 249798 197072 249854 197472
rect 254766 197072 254822 197472
rect 259734 197072 259790 197472
rect 264702 197072 264758 197472
rect 269670 197072 269726 197472
rect 274546 197072 274602 197472
rect 279514 197072 279570 197472
rect 284482 197072 284538 197472
rect 289450 197072 289506 197472
rect 294418 197072 294474 197472
rect 299294 197072 299350 197472
rect 304262 197072 304318 197472
rect 309230 197072 309286 197472
rect 314198 197072 314254 197472
rect 2410 0 2466 400
rect 7286 0 7342 400
rect 12254 0 12310 400
rect 17222 0 17278 400
rect 22190 0 22246 400
rect 27066 0 27122 400
rect 32034 0 32090 400
rect 37002 0 37058 400
rect 41970 0 42026 400
rect 46938 0 46994 400
rect 51814 0 51870 400
rect 56782 0 56838 400
rect 61750 0 61806 400
rect 66718 0 66774 400
rect 71686 0 71742 400
rect 76562 0 76618 400
rect 81530 0 81586 400
rect 86498 0 86554 400
rect 91466 0 91522 400
rect 96434 0 96490 400
rect 101310 0 101366 400
rect 106278 0 106334 400
rect 111246 0 111302 400
rect 116214 0 116270 400
rect 121182 0 121238 400
rect 126058 0 126114 400
rect 131026 0 131082 400
rect 135994 0 136050 400
rect 140962 0 141018 400
rect 145930 0 145986 400
rect 150806 0 150862 400
rect 155774 0 155830 400
rect 160742 0 160798 400
rect 165710 0 165766 400
rect 170678 0 170734 400
rect 175554 0 175610 400
rect 180522 0 180578 400
rect 185490 0 185546 400
rect 190458 0 190514 400
rect 195426 0 195482 400
rect 200302 0 200358 400
rect 205270 0 205326 400
rect 210238 0 210294 400
rect 215206 0 215262 400
rect 220174 0 220230 400
rect 225050 0 225106 400
rect 230018 0 230074 400
rect 234986 0 235042 400
rect 239954 0 240010 400
rect 244922 0 244978 400
rect 249798 0 249854 400
rect 254766 0 254822 400
rect 259734 0 259790 400
rect 264702 0 264758 400
rect 269670 0 269726 400
rect 274546 0 274602 400
rect 279514 0 279570 400
rect 284482 0 284538 400
rect 289450 0 289506 400
rect 294418 0 294474 400
rect 299294 0 299350 400
rect 304262 0 304318 400
rect 309230 0 309286 400
rect 314198 0 314254 400
<< obsm2 >>
rect 296 197016 2354 197470
rect 2522 197016 7230 197470
rect 7398 197016 12198 197470
rect 12366 197016 17166 197470
rect 17334 197016 22134 197470
rect 22302 197016 27010 197470
rect 27178 197016 31978 197470
rect 32146 197016 36946 197470
rect 37114 197016 41914 197470
rect 42082 197016 46882 197470
rect 47050 197016 51758 197470
rect 51926 197016 56726 197470
rect 56894 197016 61694 197470
rect 61862 197016 66662 197470
rect 66830 197016 71630 197470
rect 71798 197016 76506 197470
rect 76674 197016 81474 197470
rect 81642 197016 86442 197470
rect 86610 197016 91410 197470
rect 91578 197016 96378 197470
rect 96546 197016 101254 197470
rect 101422 197016 106222 197470
rect 106390 197016 111190 197470
rect 111358 197016 116158 197470
rect 116326 197016 121126 197470
rect 121294 197016 126002 197470
rect 126170 197016 130970 197470
rect 131138 197016 135938 197470
rect 136106 197016 140906 197470
rect 141074 197016 145874 197470
rect 146042 197016 150750 197470
rect 150918 197016 155718 197470
rect 155886 197016 160686 197470
rect 160854 197016 165654 197470
rect 165822 197016 170622 197470
rect 170790 197016 175498 197470
rect 175666 197016 180466 197470
rect 180634 197016 185434 197470
rect 185602 197016 190402 197470
rect 190570 197016 195370 197470
rect 195538 197016 200246 197470
rect 200414 197016 205214 197470
rect 205382 197016 210182 197470
rect 210350 197016 215150 197470
rect 215318 197016 220118 197470
rect 220286 197016 224994 197470
rect 225162 197016 229962 197470
rect 230130 197016 234930 197470
rect 235098 197016 239898 197470
rect 240066 197016 244866 197470
rect 245034 197016 249742 197470
rect 249910 197016 254710 197470
rect 254878 197016 259678 197470
rect 259846 197016 264646 197470
rect 264814 197016 269614 197470
rect 269782 197016 274490 197470
rect 274658 197016 279458 197470
rect 279626 197016 284426 197470
rect 284594 197016 289394 197470
rect 289562 197016 294362 197470
rect 294530 197016 299238 197470
rect 299406 197016 304206 197470
rect 304374 197016 309174 197470
rect 309342 197016 314142 197470
rect 314310 197016 316184 197470
rect 296 456 316184 197016
rect 296 31 2354 456
rect 2522 31 7230 456
rect 7398 31 12198 456
rect 12366 31 17166 456
rect 17334 31 22134 456
rect 22302 31 27010 456
rect 27178 31 31978 456
rect 32146 31 36946 456
rect 37114 31 41914 456
rect 42082 31 46882 456
rect 47050 31 51758 456
rect 51926 31 56726 456
rect 56894 31 61694 456
rect 61862 31 66662 456
rect 66830 31 71630 456
rect 71798 31 76506 456
rect 76674 31 81474 456
rect 81642 31 86442 456
rect 86610 31 91410 456
rect 91578 31 96378 456
rect 96546 31 101254 456
rect 101422 31 106222 456
rect 106390 31 111190 456
rect 111358 31 116158 456
rect 116326 31 121126 456
rect 121294 31 126002 456
rect 126170 31 130970 456
rect 131138 31 135938 456
rect 136106 31 140906 456
rect 141074 31 145874 456
rect 146042 31 150750 456
rect 150918 31 155718 456
rect 155886 31 160686 456
rect 160854 31 165654 456
rect 165822 31 170622 456
rect 170790 31 175498 456
rect 175666 31 180466 456
rect 180634 31 185434 456
rect 185602 31 190402 456
rect 190570 31 195370 456
rect 195538 31 200246 456
rect 200414 31 205214 456
rect 205382 31 210182 456
rect 210350 31 215150 456
rect 215318 31 220118 456
rect 220286 31 224994 456
rect 225162 31 229962 456
rect 230130 31 234930 456
rect 235098 31 239898 456
rect 240066 31 244866 456
rect 245034 31 249742 456
rect 249910 31 254710 456
rect 254878 31 259678 456
rect 259846 31 264646 456
rect 264814 31 269614 456
rect 269782 31 274490 456
rect 274658 31 279458 456
rect 279626 31 284426 456
rect 284594 31 289394 456
rect 289562 31 294362 456
rect 294530 31 299238 456
rect 299406 31 304206 456
rect 304374 31 309174 456
rect 309342 31 314142 456
rect 314310 31 316184 456
<< metal3 >>
rect 316356 191904 316756 192024
rect 316356 180888 316756 181008
rect 316356 170008 316756 170128
rect 316356 158992 316756 159112
rect 316356 147976 316756 148096
rect 316356 137096 316756 137216
rect 316356 126080 316756 126200
rect 316356 115064 316756 115184
rect 316356 104184 316756 104304
rect 0 98744 400 98864
rect 316356 93168 316756 93288
rect 316356 82152 316756 82272
rect 316356 71272 316756 71392
rect 316356 60256 316756 60376
rect 316356 49240 316756 49360
rect 316356 38360 316756 38480
rect 316356 27344 316756 27464
rect 316356 16328 316756 16448
rect 316356 5448 316756 5568
<< obsm3 >>
rect 381 192104 316356 197437
rect 381 191824 316276 192104
rect 381 181088 316356 191824
rect 381 180808 316276 181088
rect 381 170208 316356 180808
rect 381 169928 316276 170208
rect 381 159192 316356 169928
rect 381 158912 316276 159192
rect 381 148176 316356 158912
rect 381 147896 316276 148176
rect 381 137296 316356 147896
rect 381 137016 316276 137296
rect 381 126280 316356 137016
rect 381 126000 316276 126280
rect 381 115264 316356 126000
rect 381 114984 316276 115264
rect 381 104384 316356 114984
rect 381 104104 316276 104384
rect 381 98944 316356 104104
rect 480 98664 316356 98944
rect 381 93368 316356 98664
rect 381 93088 316276 93368
rect 381 82352 316356 93088
rect 381 82072 316276 82352
rect 381 71472 316356 82072
rect 381 71192 316276 71472
rect 381 60456 316356 71192
rect 381 60176 316276 60456
rect 381 49440 316356 60176
rect 381 49160 316276 49440
rect 381 38560 316356 49160
rect 381 38280 316276 38560
rect 381 27544 316356 38280
rect 381 27264 316276 27544
rect 381 16528 316356 27264
rect 381 16248 316276 16528
rect 381 5648 316356 16248
rect 381 5368 316276 5648
rect 381 35 316356 5368
<< metal4 >>
rect 4738 20080 5358 177392
rect 22738 20080 23358 177392
rect 40738 20080 41358 177392
rect 58738 20080 59358 177392
rect 76738 20080 77358 177392
rect 94738 20080 95358 177392
rect 112738 20080 113358 177392
rect 130738 20080 131358 177392
rect 148738 20080 149358 177392
rect 166738 20080 167358 177392
rect 184738 20080 185358 177392
rect 202738 20080 203358 177392
rect 220738 20080 221358 177392
rect 238738 20080 239358 177392
rect 256738 20080 257358 177392
rect 274738 20080 275358 177392
rect 292738 20080 293358 177392
rect 310738 20080 311358 177392
<< obsm4 >>
rect 2635 177472 313845 197437
rect 2635 20000 4658 177472
rect 5438 20000 22658 177472
rect 23438 20000 40658 177472
rect 41438 20000 58658 177472
rect 59438 20000 76658 177472
rect 77438 20000 94658 177472
rect 95438 20000 112658 177472
rect 113438 20000 130658 177472
rect 131438 20000 148658 177472
rect 149438 20000 166658 177472
rect 167438 20000 184658 177472
rect 185438 20000 202658 177472
rect 203438 20000 220658 177472
rect 221438 20000 238658 177472
rect 239438 20000 256658 177472
rect 257438 20000 274658 177472
rect 275438 20000 292658 177472
rect 293438 20000 310658 177472
rect 311438 20000 313845 177472
rect 2635 171 313845 20000
<< labels >>
rlabel metal3 s 316356 104184 316756 104304 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 316356 115064 316756 115184 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 316356 126080 316756 126200 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 316356 137096 316756 137216 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 316356 147976 316756 148096 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 316356 158992 316756 159112 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 316356 170008 316756 170128 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 316356 180888 316756 181008 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 316356 191904 316756 192024 6 A0[8]
port 9 nsew signal input
rlabel metal3 s 0 98744 400 98864 6 CLK
port 10 nsew signal input
rlabel metal2 s 2410 0 2466 400 6 Di0[0]
port 11 nsew signal input
rlabel metal2 s 51814 0 51870 400 6 Di0[10]
port 12 nsew signal input
rlabel metal2 s 56782 0 56838 400 6 Di0[11]
port 13 nsew signal input
rlabel metal2 s 61750 0 61806 400 6 Di0[12]
port 14 nsew signal input
rlabel metal2 s 66718 0 66774 400 6 Di0[13]
port 15 nsew signal input
rlabel metal2 s 71686 0 71742 400 6 Di0[14]
port 16 nsew signal input
rlabel metal2 s 76562 0 76618 400 6 Di0[15]
port 17 nsew signal input
rlabel metal2 s 81530 0 81586 400 6 Di0[16]
port 18 nsew signal input
rlabel metal2 s 86498 0 86554 400 6 Di0[17]
port 19 nsew signal input
rlabel metal2 s 91466 0 91522 400 6 Di0[18]
port 20 nsew signal input
rlabel metal2 s 96434 0 96490 400 6 Di0[19]
port 21 nsew signal input
rlabel metal2 s 7286 0 7342 400 6 Di0[1]
port 22 nsew signal input
rlabel metal2 s 101310 0 101366 400 6 Di0[20]
port 23 nsew signal input
rlabel metal2 s 106278 0 106334 400 6 Di0[21]
port 24 nsew signal input
rlabel metal2 s 111246 0 111302 400 6 Di0[22]
port 25 nsew signal input
rlabel metal2 s 116214 0 116270 400 6 Di0[23]
port 26 nsew signal input
rlabel metal2 s 121182 0 121238 400 6 Di0[24]
port 27 nsew signal input
rlabel metal2 s 126058 0 126114 400 6 Di0[25]
port 28 nsew signal input
rlabel metal2 s 131026 0 131082 400 6 Di0[26]
port 29 nsew signal input
rlabel metal2 s 135994 0 136050 400 6 Di0[27]
port 30 nsew signal input
rlabel metal2 s 140962 0 141018 400 6 Di0[28]
port 31 nsew signal input
rlabel metal2 s 145930 0 145986 400 6 Di0[29]
port 32 nsew signal input
rlabel metal2 s 12254 0 12310 400 6 Di0[2]
port 33 nsew signal input
rlabel metal2 s 150806 0 150862 400 6 Di0[30]
port 34 nsew signal input
rlabel metal2 s 155774 0 155830 400 6 Di0[31]
port 35 nsew signal input
rlabel metal2 s 160742 0 160798 400 6 Di0[32]
port 36 nsew signal input
rlabel metal2 s 165710 0 165766 400 6 Di0[33]
port 37 nsew signal input
rlabel metal2 s 170678 0 170734 400 6 Di0[34]
port 38 nsew signal input
rlabel metal2 s 175554 0 175610 400 6 Di0[35]
port 39 nsew signal input
rlabel metal2 s 180522 0 180578 400 6 Di0[36]
port 40 nsew signal input
rlabel metal2 s 185490 0 185546 400 6 Di0[37]
port 41 nsew signal input
rlabel metal2 s 190458 0 190514 400 6 Di0[38]
port 42 nsew signal input
rlabel metal2 s 195426 0 195482 400 6 Di0[39]
port 43 nsew signal input
rlabel metal2 s 17222 0 17278 400 6 Di0[3]
port 44 nsew signal input
rlabel metal2 s 200302 0 200358 400 6 Di0[40]
port 45 nsew signal input
rlabel metal2 s 205270 0 205326 400 6 Di0[41]
port 46 nsew signal input
rlabel metal2 s 210238 0 210294 400 6 Di0[42]
port 47 nsew signal input
rlabel metal2 s 215206 0 215262 400 6 Di0[43]
port 48 nsew signal input
rlabel metal2 s 220174 0 220230 400 6 Di0[44]
port 49 nsew signal input
rlabel metal2 s 225050 0 225106 400 6 Di0[45]
port 50 nsew signal input
rlabel metal2 s 230018 0 230074 400 6 Di0[46]
port 51 nsew signal input
rlabel metal2 s 234986 0 235042 400 6 Di0[47]
port 52 nsew signal input
rlabel metal2 s 239954 0 240010 400 6 Di0[48]
port 53 nsew signal input
rlabel metal2 s 244922 0 244978 400 6 Di0[49]
port 54 nsew signal input
rlabel metal2 s 22190 0 22246 400 6 Di0[4]
port 55 nsew signal input
rlabel metal2 s 249798 0 249854 400 6 Di0[50]
port 56 nsew signal input
rlabel metal2 s 254766 0 254822 400 6 Di0[51]
port 57 nsew signal input
rlabel metal2 s 259734 0 259790 400 6 Di0[52]
port 58 nsew signal input
rlabel metal2 s 264702 0 264758 400 6 Di0[53]
port 59 nsew signal input
rlabel metal2 s 269670 0 269726 400 6 Di0[54]
port 60 nsew signal input
rlabel metal2 s 274546 0 274602 400 6 Di0[55]
port 61 nsew signal input
rlabel metal2 s 279514 0 279570 400 6 Di0[56]
port 62 nsew signal input
rlabel metal2 s 284482 0 284538 400 6 Di0[57]
port 63 nsew signal input
rlabel metal2 s 289450 0 289506 400 6 Di0[58]
port 64 nsew signal input
rlabel metal2 s 294418 0 294474 400 6 Di0[59]
port 65 nsew signal input
rlabel metal2 s 27066 0 27122 400 6 Di0[5]
port 66 nsew signal input
rlabel metal2 s 299294 0 299350 400 6 Di0[60]
port 67 nsew signal input
rlabel metal2 s 304262 0 304318 400 6 Di0[61]
port 68 nsew signal input
rlabel metal2 s 309230 0 309286 400 6 Di0[62]
port 69 nsew signal input
rlabel metal2 s 314198 0 314254 400 6 Di0[63]
port 70 nsew signal input
rlabel metal2 s 32034 0 32090 400 6 Di0[6]
port 71 nsew signal input
rlabel metal2 s 37002 0 37058 400 6 Di0[7]
port 72 nsew signal input
rlabel metal2 s 41970 0 42026 400 6 Di0[8]
port 73 nsew signal input
rlabel metal2 s 46938 0 46994 400 6 Di0[9]
port 74 nsew signal input
rlabel metal2 s 2410 197072 2466 197472 6 Do0[0]
port 75 nsew signal output
rlabel metal2 s 51814 197072 51870 197472 6 Do0[10]
port 76 nsew signal output
rlabel metal2 s 56782 197072 56838 197472 6 Do0[11]
port 77 nsew signal output
rlabel metal2 s 61750 197072 61806 197472 6 Do0[12]
port 78 nsew signal output
rlabel metal2 s 66718 197072 66774 197472 6 Do0[13]
port 79 nsew signal output
rlabel metal2 s 71686 197072 71742 197472 6 Do0[14]
port 80 nsew signal output
rlabel metal2 s 76562 197072 76618 197472 6 Do0[15]
port 81 nsew signal output
rlabel metal2 s 81530 197072 81586 197472 6 Do0[16]
port 82 nsew signal output
rlabel metal2 s 86498 197072 86554 197472 6 Do0[17]
port 83 nsew signal output
rlabel metal2 s 91466 197072 91522 197472 6 Do0[18]
port 84 nsew signal output
rlabel metal2 s 96434 197072 96490 197472 6 Do0[19]
port 85 nsew signal output
rlabel metal2 s 7286 197072 7342 197472 6 Do0[1]
port 86 nsew signal output
rlabel metal2 s 101310 197072 101366 197472 6 Do0[20]
port 87 nsew signal output
rlabel metal2 s 106278 197072 106334 197472 6 Do0[21]
port 88 nsew signal output
rlabel metal2 s 111246 197072 111302 197472 6 Do0[22]
port 89 nsew signal output
rlabel metal2 s 116214 197072 116270 197472 6 Do0[23]
port 90 nsew signal output
rlabel metal2 s 121182 197072 121238 197472 6 Do0[24]
port 91 nsew signal output
rlabel metal2 s 126058 197072 126114 197472 6 Do0[25]
port 92 nsew signal output
rlabel metal2 s 131026 197072 131082 197472 6 Do0[26]
port 93 nsew signal output
rlabel metal2 s 135994 197072 136050 197472 6 Do0[27]
port 94 nsew signal output
rlabel metal2 s 140962 197072 141018 197472 6 Do0[28]
port 95 nsew signal output
rlabel metal2 s 145930 197072 145986 197472 6 Do0[29]
port 96 nsew signal output
rlabel metal2 s 12254 197072 12310 197472 6 Do0[2]
port 97 nsew signal output
rlabel metal2 s 150806 197072 150862 197472 6 Do0[30]
port 98 nsew signal output
rlabel metal2 s 155774 197072 155830 197472 6 Do0[31]
port 99 nsew signal output
rlabel metal2 s 160742 197072 160798 197472 6 Do0[32]
port 100 nsew signal output
rlabel metal2 s 165710 197072 165766 197472 6 Do0[33]
port 101 nsew signal output
rlabel metal2 s 170678 197072 170734 197472 6 Do0[34]
port 102 nsew signal output
rlabel metal2 s 175554 197072 175610 197472 6 Do0[35]
port 103 nsew signal output
rlabel metal2 s 180522 197072 180578 197472 6 Do0[36]
port 104 nsew signal output
rlabel metal2 s 185490 197072 185546 197472 6 Do0[37]
port 105 nsew signal output
rlabel metal2 s 190458 197072 190514 197472 6 Do0[38]
port 106 nsew signal output
rlabel metal2 s 195426 197072 195482 197472 6 Do0[39]
port 107 nsew signal output
rlabel metal2 s 17222 197072 17278 197472 6 Do0[3]
port 108 nsew signal output
rlabel metal2 s 200302 197072 200358 197472 6 Do0[40]
port 109 nsew signal output
rlabel metal2 s 205270 197072 205326 197472 6 Do0[41]
port 110 nsew signal output
rlabel metal2 s 210238 197072 210294 197472 6 Do0[42]
port 111 nsew signal output
rlabel metal2 s 215206 197072 215262 197472 6 Do0[43]
port 112 nsew signal output
rlabel metal2 s 220174 197072 220230 197472 6 Do0[44]
port 113 nsew signal output
rlabel metal2 s 225050 197072 225106 197472 6 Do0[45]
port 114 nsew signal output
rlabel metal2 s 230018 197072 230074 197472 6 Do0[46]
port 115 nsew signal output
rlabel metal2 s 234986 197072 235042 197472 6 Do0[47]
port 116 nsew signal output
rlabel metal2 s 239954 197072 240010 197472 6 Do0[48]
port 117 nsew signal output
rlabel metal2 s 244922 197072 244978 197472 6 Do0[49]
port 118 nsew signal output
rlabel metal2 s 22190 197072 22246 197472 6 Do0[4]
port 119 nsew signal output
rlabel metal2 s 249798 197072 249854 197472 6 Do0[50]
port 120 nsew signal output
rlabel metal2 s 254766 197072 254822 197472 6 Do0[51]
port 121 nsew signal output
rlabel metal2 s 259734 197072 259790 197472 6 Do0[52]
port 122 nsew signal output
rlabel metal2 s 264702 197072 264758 197472 6 Do0[53]
port 123 nsew signal output
rlabel metal2 s 269670 197072 269726 197472 6 Do0[54]
port 124 nsew signal output
rlabel metal2 s 274546 197072 274602 197472 6 Do0[55]
port 125 nsew signal output
rlabel metal2 s 279514 197072 279570 197472 6 Do0[56]
port 126 nsew signal output
rlabel metal2 s 284482 197072 284538 197472 6 Do0[57]
port 127 nsew signal output
rlabel metal2 s 289450 197072 289506 197472 6 Do0[58]
port 128 nsew signal output
rlabel metal2 s 294418 197072 294474 197472 6 Do0[59]
port 129 nsew signal output
rlabel metal2 s 27066 197072 27122 197472 6 Do0[5]
port 130 nsew signal output
rlabel metal2 s 299294 197072 299350 197472 6 Do0[60]
port 131 nsew signal output
rlabel metal2 s 304262 197072 304318 197472 6 Do0[61]
port 132 nsew signal output
rlabel metal2 s 309230 197072 309286 197472 6 Do0[62]
port 133 nsew signal output
rlabel metal2 s 314198 197072 314254 197472 6 Do0[63]
port 134 nsew signal output
rlabel metal2 s 32034 197072 32090 197472 6 Do0[6]
port 135 nsew signal output
rlabel metal2 s 37002 197072 37058 197472 6 Do0[7]
port 136 nsew signal output
rlabel metal2 s 41970 197072 42026 197472 6 Do0[8]
port 137 nsew signal output
rlabel metal2 s 46938 197072 46994 197472 6 Do0[9]
port 138 nsew signal output
rlabel metal3 s 316356 5448 316756 5568 6 EN0
port 139 nsew signal input
rlabel metal4 s 22738 20080 23358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 58738 20080 59358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 94738 20080 95358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 130738 20080 131358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 166738 20080 167358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 202738 20080 203358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 238738 20080 239358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 274738 20080 275358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 310738 20080 311358 177392 6 VGND
port 140 nsew ground bidirectional
rlabel metal4 s 4738 20080 5358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 40738 20080 41358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 76738 20080 77358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 112738 20080 113358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 148738 20080 149358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 184738 20080 185358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 220738 20080 221358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 256738 20080 257358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal4 s 292738 20080 293358 177392 6 VPWR
port 141 nsew power bidirectional
rlabel metal3 s 316356 16328 316756 16448 6 WE0[0]
port 142 nsew signal input
rlabel metal3 s 316356 27344 316756 27464 6 WE0[1]
port 143 nsew signal input
rlabel metal3 s 316356 38360 316756 38480 6 WE0[2]
port 144 nsew signal input
rlabel metal3 s 316356 49240 316756 49360 6 WE0[3]
port 145 nsew signal input
rlabel metal3 s 316356 60256 316756 60376 6 WE0[4]
port 146 nsew signal input
rlabel metal3 s 316356 71272 316756 71392 6 WE0[5]
port 147 nsew signal input
rlabel metal3 s 316356 82152 316756 82272 6 WE0[6]
port 148 nsew signal input
rlabel metal3 s 316356 93168 316756 93288 6 WE0[7]
port 149 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 316756 197472
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 190679036
string GDS_FILE /mnt/dffram/build/512x64_DEFAULT/openlane/runs/RUN_2022.06.07_03.41.15/results/signoff/RAM512.magic.gds
string GDS_START 165654
<< end >>

