magic
tech sky130A
magscale 1 2
timestamp 1654573573
<< obsli1 >>
rect 1104 2159 118864 117521
<< obsm1 >>
rect 474 1572 119678 117552
<< metal2 >>
rect 478 119200 534 120000
rect 1398 119200 1454 120000
rect 2318 119200 2374 120000
rect 3238 119200 3294 120000
rect 4158 119200 4214 120000
rect 5078 119200 5134 120000
rect 5998 119200 6054 120000
rect 6918 119200 6974 120000
rect 7838 119200 7894 120000
rect 8758 119200 8814 120000
rect 9678 119200 9734 120000
rect 10598 119200 10654 120000
rect 11518 119200 11574 120000
rect 12438 119200 12494 120000
rect 13358 119200 13414 120000
rect 14278 119200 14334 120000
rect 15198 119200 15254 120000
rect 16118 119200 16174 120000
rect 17038 119200 17094 120000
rect 17958 119200 18014 120000
rect 18878 119200 18934 120000
rect 19798 119200 19854 120000
rect 20718 119200 20774 120000
rect 21638 119200 21694 120000
rect 22558 119200 22614 120000
rect 23478 119200 23534 120000
rect 24398 119200 24454 120000
rect 25318 119200 25374 120000
rect 26238 119200 26294 120000
rect 27158 119200 27214 120000
rect 28078 119200 28134 120000
rect 28998 119200 29054 120000
rect 29918 119200 29974 120000
rect 30930 119200 30986 120000
rect 31850 119200 31906 120000
rect 32770 119200 32826 120000
rect 33690 119200 33746 120000
rect 34610 119200 34666 120000
rect 35530 119200 35586 120000
rect 36450 119200 36506 120000
rect 37370 119200 37426 120000
rect 38290 119200 38346 120000
rect 39210 119200 39266 120000
rect 40130 119200 40186 120000
rect 41050 119200 41106 120000
rect 41970 119200 42026 120000
rect 42890 119200 42946 120000
rect 43810 119200 43866 120000
rect 44730 119200 44786 120000
rect 45650 119200 45706 120000
rect 46570 119200 46626 120000
rect 47490 119200 47546 120000
rect 48410 119200 48466 120000
rect 49330 119200 49386 120000
rect 50250 119200 50306 120000
rect 51170 119200 51226 120000
rect 52090 119200 52146 120000
rect 53010 119200 53066 120000
rect 53930 119200 53986 120000
rect 54850 119200 54906 120000
rect 55770 119200 55826 120000
rect 56690 119200 56746 120000
rect 57610 119200 57666 120000
rect 58530 119200 58586 120000
rect 59450 119200 59506 120000
rect 60462 119200 60518 120000
rect 61382 119200 61438 120000
rect 62302 119200 62358 120000
rect 63222 119200 63278 120000
rect 64142 119200 64198 120000
rect 65062 119200 65118 120000
rect 65982 119200 66038 120000
rect 66902 119200 66958 120000
rect 67822 119200 67878 120000
rect 68742 119200 68798 120000
rect 69662 119200 69718 120000
rect 70582 119200 70638 120000
rect 71502 119200 71558 120000
rect 72422 119200 72478 120000
rect 73342 119200 73398 120000
rect 74262 119200 74318 120000
rect 75182 119200 75238 120000
rect 76102 119200 76158 120000
rect 77022 119200 77078 120000
rect 77942 119200 77998 120000
rect 78862 119200 78918 120000
rect 79782 119200 79838 120000
rect 80702 119200 80758 120000
rect 81622 119200 81678 120000
rect 82542 119200 82598 120000
rect 83462 119200 83518 120000
rect 84382 119200 84438 120000
rect 85302 119200 85358 120000
rect 86222 119200 86278 120000
rect 87142 119200 87198 120000
rect 88062 119200 88118 120000
rect 88982 119200 89038 120000
rect 89902 119200 89958 120000
rect 90914 119200 90970 120000
rect 91834 119200 91890 120000
rect 92754 119200 92810 120000
rect 93674 119200 93730 120000
rect 94594 119200 94650 120000
rect 95514 119200 95570 120000
rect 96434 119200 96490 120000
rect 97354 119200 97410 120000
rect 98274 119200 98330 120000
rect 99194 119200 99250 120000
rect 100114 119200 100170 120000
rect 101034 119200 101090 120000
rect 101954 119200 102010 120000
rect 102874 119200 102930 120000
rect 103794 119200 103850 120000
rect 104714 119200 104770 120000
rect 105634 119200 105690 120000
rect 106554 119200 106610 120000
rect 107474 119200 107530 120000
rect 108394 119200 108450 120000
rect 109314 119200 109370 120000
rect 110234 119200 110290 120000
rect 111154 119200 111210 120000
rect 112074 119200 112130 120000
rect 112994 119200 113050 120000
rect 113914 119200 113970 120000
rect 114834 119200 114890 120000
rect 115754 119200 115810 120000
rect 116674 119200 116730 120000
rect 117594 119200 117650 120000
rect 118514 119200 118570 120000
rect 119434 119200 119490 120000
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 5078 0 5134 800
rect 6090 0 6146 800
rect 7010 0 7066 800
rect 7930 0 7986 800
rect 8850 0 8906 800
rect 9770 0 9826 800
rect 10782 0 10838 800
rect 11702 0 11758 800
rect 12622 0 12678 800
rect 13542 0 13598 800
rect 14462 0 14518 800
rect 15474 0 15530 800
rect 16394 0 16450 800
rect 17314 0 17370 800
rect 18234 0 18290 800
rect 19154 0 19210 800
rect 20074 0 20130 800
rect 21086 0 21142 800
rect 22006 0 22062 800
rect 22926 0 22982 800
rect 23846 0 23902 800
rect 24766 0 24822 800
rect 25778 0 25834 800
rect 26698 0 26754 800
rect 27618 0 27674 800
rect 28538 0 28594 800
rect 29458 0 29514 800
rect 30470 0 30526 800
rect 31390 0 31446 800
rect 32310 0 32366 800
rect 33230 0 33286 800
rect 34150 0 34206 800
rect 35070 0 35126 800
rect 36082 0 36138 800
rect 37002 0 37058 800
rect 37922 0 37978 800
rect 38842 0 38898 800
rect 39762 0 39818 800
rect 40774 0 40830 800
rect 41694 0 41750 800
rect 42614 0 42670 800
rect 43534 0 43590 800
rect 44454 0 44510 800
rect 45466 0 45522 800
rect 46386 0 46442 800
rect 47306 0 47362 800
rect 48226 0 48282 800
rect 49146 0 49202 800
rect 50066 0 50122 800
rect 51078 0 51134 800
rect 51998 0 52054 800
rect 52918 0 52974 800
rect 53838 0 53894 800
rect 54758 0 54814 800
rect 55770 0 55826 800
rect 56690 0 56746 800
rect 57610 0 57666 800
rect 58530 0 58586 800
rect 59450 0 59506 800
rect 60462 0 60518 800
rect 61382 0 61438 800
rect 62302 0 62358 800
rect 63222 0 63278 800
rect 64142 0 64198 800
rect 65062 0 65118 800
rect 66074 0 66130 800
rect 66994 0 67050 800
rect 67914 0 67970 800
rect 68834 0 68890 800
rect 69754 0 69810 800
rect 70766 0 70822 800
rect 71686 0 71742 800
rect 72606 0 72662 800
rect 73526 0 73582 800
rect 74446 0 74502 800
rect 75458 0 75514 800
rect 76378 0 76434 800
rect 77298 0 77354 800
rect 78218 0 78274 800
rect 79138 0 79194 800
rect 80058 0 80114 800
rect 81070 0 81126 800
rect 81990 0 82046 800
rect 82910 0 82966 800
rect 83830 0 83886 800
rect 84750 0 84806 800
rect 85762 0 85818 800
rect 86682 0 86738 800
rect 87602 0 87658 800
rect 88522 0 88578 800
rect 89442 0 89498 800
rect 90454 0 90510 800
rect 91374 0 91430 800
rect 92294 0 92350 800
rect 93214 0 93270 800
rect 94134 0 94190 800
rect 95054 0 95110 800
rect 96066 0 96122 800
rect 96986 0 97042 800
rect 97906 0 97962 800
rect 98826 0 98882 800
rect 99746 0 99802 800
rect 100758 0 100814 800
rect 101678 0 101734 800
rect 102598 0 102654 800
rect 103518 0 103574 800
rect 104438 0 104494 800
rect 105450 0 105506 800
rect 106370 0 106426 800
rect 107290 0 107346 800
rect 108210 0 108266 800
rect 109130 0 109186 800
rect 110050 0 110106 800
rect 111062 0 111118 800
rect 111982 0 112038 800
rect 112902 0 112958 800
rect 113822 0 113878 800
rect 114742 0 114798 800
rect 115754 0 115810 800
rect 116674 0 116730 800
rect 117594 0 117650 800
rect 118514 0 118570 800
rect 119434 0 119490 800
<< obsm2 >>
rect 590 119144 1342 119513
rect 1510 119144 2262 119513
rect 2430 119144 3182 119513
rect 3350 119144 4102 119513
rect 4270 119144 5022 119513
rect 5190 119144 5942 119513
rect 6110 119144 6862 119513
rect 7030 119144 7782 119513
rect 7950 119144 8702 119513
rect 8870 119144 9622 119513
rect 9790 119144 10542 119513
rect 10710 119144 11462 119513
rect 11630 119144 12382 119513
rect 12550 119144 13302 119513
rect 13470 119144 14222 119513
rect 14390 119144 15142 119513
rect 15310 119144 16062 119513
rect 16230 119144 16982 119513
rect 17150 119144 17902 119513
rect 18070 119144 18822 119513
rect 18990 119144 19742 119513
rect 19910 119144 20662 119513
rect 20830 119144 21582 119513
rect 21750 119144 22502 119513
rect 22670 119144 23422 119513
rect 23590 119144 24342 119513
rect 24510 119144 25262 119513
rect 25430 119144 26182 119513
rect 26350 119144 27102 119513
rect 27270 119144 28022 119513
rect 28190 119144 28942 119513
rect 29110 119144 29862 119513
rect 30030 119144 30874 119513
rect 31042 119144 31794 119513
rect 31962 119144 32714 119513
rect 32882 119144 33634 119513
rect 33802 119144 34554 119513
rect 34722 119144 35474 119513
rect 35642 119144 36394 119513
rect 36562 119144 37314 119513
rect 37482 119144 38234 119513
rect 38402 119144 39154 119513
rect 39322 119144 40074 119513
rect 40242 119144 40994 119513
rect 41162 119144 41914 119513
rect 42082 119144 42834 119513
rect 43002 119144 43754 119513
rect 43922 119144 44674 119513
rect 44842 119144 45594 119513
rect 45762 119144 46514 119513
rect 46682 119144 47434 119513
rect 47602 119144 48354 119513
rect 48522 119144 49274 119513
rect 49442 119144 50194 119513
rect 50362 119144 51114 119513
rect 51282 119144 52034 119513
rect 52202 119144 52954 119513
rect 53122 119144 53874 119513
rect 54042 119144 54794 119513
rect 54962 119144 55714 119513
rect 55882 119144 56634 119513
rect 56802 119144 57554 119513
rect 57722 119144 58474 119513
rect 58642 119144 59394 119513
rect 59562 119144 60406 119513
rect 60574 119144 61326 119513
rect 61494 119144 62246 119513
rect 62414 119144 63166 119513
rect 63334 119144 64086 119513
rect 64254 119144 65006 119513
rect 65174 119144 65926 119513
rect 66094 119144 66846 119513
rect 67014 119144 67766 119513
rect 67934 119144 68686 119513
rect 68854 119144 69606 119513
rect 69774 119144 70526 119513
rect 70694 119144 71446 119513
rect 71614 119144 72366 119513
rect 72534 119144 73286 119513
rect 73454 119144 74206 119513
rect 74374 119144 75126 119513
rect 75294 119144 76046 119513
rect 76214 119144 76966 119513
rect 77134 119144 77886 119513
rect 78054 119144 78806 119513
rect 78974 119144 79726 119513
rect 79894 119144 80646 119513
rect 80814 119144 81566 119513
rect 81734 119144 82486 119513
rect 82654 119144 83406 119513
rect 83574 119144 84326 119513
rect 84494 119144 85246 119513
rect 85414 119144 86166 119513
rect 86334 119144 87086 119513
rect 87254 119144 88006 119513
rect 88174 119144 88926 119513
rect 89094 119144 89846 119513
rect 90014 119144 90858 119513
rect 91026 119144 91778 119513
rect 91946 119144 92698 119513
rect 92866 119144 93618 119513
rect 93786 119144 94538 119513
rect 94706 119144 95458 119513
rect 95626 119144 96378 119513
rect 96546 119144 97298 119513
rect 97466 119144 98218 119513
rect 98386 119144 99138 119513
rect 99306 119144 100058 119513
rect 100226 119144 100978 119513
rect 101146 119144 101898 119513
rect 102066 119144 102818 119513
rect 102986 119144 103738 119513
rect 103906 119144 104658 119513
rect 104826 119144 105578 119513
rect 105746 119144 106498 119513
rect 106666 119144 107418 119513
rect 107586 119144 108338 119513
rect 108506 119144 109258 119513
rect 109426 119144 110178 119513
rect 110346 119144 111098 119513
rect 111266 119144 112018 119513
rect 112186 119144 112938 119513
rect 113106 119144 113858 119513
rect 114026 119144 114778 119513
rect 114946 119144 115698 119513
rect 115866 119144 116618 119513
rect 116786 119144 117538 119513
rect 117706 119144 118458 119513
rect 118626 119144 119378 119513
rect 119546 119144 119672 119513
rect 480 856 119672 119144
rect 590 734 1342 856
rect 1510 734 2262 856
rect 2430 734 3182 856
rect 3350 734 4102 856
rect 4270 734 5022 856
rect 5190 734 6034 856
rect 6202 734 6954 856
rect 7122 734 7874 856
rect 8042 734 8794 856
rect 8962 734 9714 856
rect 9882 734 10726 856
rect 10894 734 11646 856
rect 11814 734 12566 856
rect 12734 734 13486 856
rect 13654 734 14406 856
rect 14574 734 15418 856
rect 15586 734 16338 856
rect 16506 734 17258 856
rect 17426 734 18178 856
rect 18346 734 19098 856
rect 19266 734 20018 856
rect 20186 734 21030 856
rect 21198 734 21950 856
rect 22118 734 22870 856
rect 23038 734 23790 856
rect 23958 734 24710 856
rect 24878 734 25722 856
rect 25890 734 26642 856
rect 26810 734 27562 856
rect 27730 734 28482 856
rect 28650 734 29402 856
rect 29570 734 30414 856
rect 30582 734 31334 856
rect 31502 734 32254 856
rect 32422 734 33174 856
rect 33342 734 34094 856
rect 34262 734 35014 856
rect 35182 734 36026 856
rect 36194 734 36946 856
rect 37114 734 37866 856
rect 38034 734 38786 856
rect 38954 734 39706 856
rect 39874 734 40718 856
rect 40886 734 41638 856
rect 41806 734 42558 856
rect 42726 734 43478 856
rect 43646 734 44398 856
rect 44566 734 45410 856
rect 45578 734 46330 856
rect 46498 734 47250 856
rect 47418 734 48170 856
rect 48338 734 49090 856
rect 49258 734 50010 856
rect 50178 734 51022 856
rect 51190 734 51942 856
rect 52110 734 52862 856
rect 53030 734 53782 856
rect 53950 734 54702 856
rect 54870 734 55714 856
rect 55882 734 56634 856
rect 56802 734 57554 856
rect 57722 734 58474 856
rect 58642 734 59394 856
rect 59562 734 60406 856
rect 60574 734 61326 856
rect 61494 734 62246 856
rect 62414 734 63166 856
rect 63334 734 64086 856
rect 64254 734 65006 856
rect 65174 734 66018 856
rect 66186 734 66938 856
rect 67106 734 67858 856
rect 68026 734 68778 856
rect 68946 734 69698 856
rect 69866 734 70710 856
rect 70878 734 71630 856
rect 71798 734 72550 856
rect 72718 734 73470 856
rect 73638 734 74390 856
rect 74558 734 75402 856
rect 75570 734 76322 856
rect 76490 734 77242 856
rect 77410 734 78162 856
rect 78330 734 79082 856
rect 79250 734 80002 856
rect 80170 734 81014 856
rect 81182 734 81934 856
rect 82102 734 82854 856
rect 83022 734 83774 856
rect 83942 734 84694 856
rect 84862 734 85706 856
rect 85874 734 86626 856
rect 86794 734 87546 856
rect 87714 734 88466 856
rect 88634 734 89386 856
rect 89554 734 90398 856
rect 90566 734 91318 856
rect 91486 734 92238 856
rect 92406 734 93158 856
rect 93326 734 94078 856
rect 94246 734 94998 856
rect 95166 734 96010 856
rect 96178 734 96930 856
rect 97098 734 97850 856
rect 98018 734 98770 856
rect 98938 734 99690 856
rect 99858 734 100702 856
rect 100870 734 101622 856
rect 101790 734 102542 856
rect 102710 734 103462 856
rect 103630 734 104382 856
rect 104550 734 105394 856
rect 105562 734 106314 856
rect 106482 734 107234 856
rect 107402 734 108154 856
rect 108322 734 109074 856
rect 109242 734 109994 856
rect 110162 734 111006 856
rect 111174 734 111926 856
rect 112094 734 112846 856
rect 113014 734 113766 856
rect 113934 734 114686 856
rect 114854 734 115698 856
rect 115866 734 116618 856
rect 116786 734 117538 856
rect 117706 734 118458 856
rect 118626 734 119378 856
rect 119546 734 119672 856
<< metal3 >>
rect 119200 119416 120000 119536
rect 119200 118464 120000 118584
rect 119200 117512 120000 117632
rect 119200 116560 120000 116680
rect 119200 115608 120000 115728
rect 119200 114656 120000 114776
rect 119200 113704 120000 113824
rect 119200 112752 120000 112872
rect 119200 111800 120000 111920
rect 119200 110984 120000 111104
rect 119200 110032 120000 110152
rect 119200 109080 120000 109200
rect 119200 108128 120000 108248
rect 119200 107176 120000 107296
rect 119200 106224 120000 106344
rect 119200 105272 120000 105392
rect 119200 104320 120000 104440
rect 119200 103368 120000 103488
rect 119200 102552 120000 102672
rect 119200 101600 120000 101720
rect 119200 100648 120000 100768
rect 119200 99696 120000 99816
rect 119200 98744 120000 98864
rect 119200 97792 120000 97912
rect 119200 96840 120000 96960
rect 119200 95888 120000 96008
rect 119200 94936 120000 95056
rect 119200 94120 120000 94240
rect 119200 93168 120000 93288
rect 119200 92216 120000 92336
rect 119200 91264 120000 91384
rect 119200 90312 120000 90432
rect 119200 89360 120000 89480
rect 119200 88408 120000 88528
rect 119200 87456 120000 87576
rect 119200 86504 120000 86624
rect 119200 85688 120000 85808
rect 119200 84736 120000 84856
rect 119200 83784 120000 83904
rect 119200 82832 120000 82952
rect 119200 81880 120000 82000
rect 119200 80928 120000 81048
rect 119200 79976 120000 80096
rect 119200 79024 120000 79144
rect 119200 78072 120000 78192
rect 119200 77256 120000 77376
rect 119200 76304 120000 76424
rect 119200 75352 120000 75472
rect 119200 74400 120000 74520
rect 119200 73448 120000 73568
rect 119200 72496 120000 72616
rect 119200 71544 120000 71664
rect 119200 70592 120000 70712
rect 119200 69640 120000 69760
rect 119200 68824 120000 68944
rect 119200 67872 120000 67992
rect 119200 66920 120000 67040
rect 119200 65968 120000 66088
rect 119200 65016 120000 65136
rect 119200 64064 120000 64184
rect 119200 63112 120000 63232
rect 119200 62160 120000 62280
rect 119200 61208 120000 61328
rect 119200 60392 120000 60512
rect 119200 59440 120000 59560
rect 119200 58488 120000 58608
rect 119200 57536 120000 57656
rect 119200 56584 120000 56704
rect 119200 55632 120000 55752
rect 119200 54680 120000 54800
rect 119200 53728 120000 53848
rect 119200 52776 120000 52896
rect 119200 51824 120000 51944
rect 119200 51008 120000 51128
rect 119200 50056 120000 50176
rect 119200 49104 120000 49224
rect 119200 48152 120000 48272
rect 119200 47200 120000 47320
rect 119200 46248 120000 46368
rect 119200 45296 120000 45416
rect 119200 44344 120000 44464
rect 119200 43392 120000 43512
rect 119200 42576 120000 42696
rect 119200 41624 120000 41744
rect 119200 40672 120000 40792
rect 119200 39720 120000 39840
rect 119200 38768 120000 38888
rect 119200 37816 120000 37936
rect 119200 36864 120000 36984
rect 119200 35912 120000 36032
rect 119200 34960 120000 35080
rect 119200 34144 120000 34264
rect 119200 33192 120000 33312
rect 119200 32240 120000 32360
rect 119200 31288 120000 31408
rect 119200 30336 120000 30456
rect 119200 29384 120000 29504
rect 119200 28432 120000 28552
rect 119200 27480 120000 27600
rect 119200 26528 120000 26648
rect 119200 25712 120000 25832
rect 119200 24760 120000 24880
rect 119200 23808 120000 23928
rect 119200 22856 120000 22976
rect 119200 21904 120000 22024
rect 119200 20952 120000 21072
rect 119200 20000 120000 20120
rect 119200 19048 120000 19168
rect 119200 18096 120000 18216
rect 119200 17280 120000 17400
rect 119200 16328 120000 16448
rect 119200 15376 120000 15496
rect 119200 14424 120000 14544
rect 119200 13472 120000 13592
rect 119200 12520 120000 12640
rect 119200 11568 120000 11688
rect 119200 10616 120000 10736
rect 119200 9664 120000 9784
rect 119200 8848 120000 8968
rect 119200 7896 120000 8016
rect 119200 6944 120000 7064
rect 119200 5992 120000 6112
rect 119200 5040 120000 5160
rect 119200 4088 120000 4208
rect 119200 3136 120000 3256
rect 119200 2184 120000 2304
rect 119200 1232 120000 1352
rect 119200 416 120000 536
<< obsm3 >>
rect 1025 119336 119120 119509
rect 1025 118664 119200 119336
rect 1025 118384 119120 118664
rect 1025 117712 119200 118384
rect 1025 117432 119120 117712
rect 1025 116760 119200 117432
rect 1025 116480 119120 116760
rect 1025 115808 119200 116480
rect 1025 115528 119120 115808
rect 1025 114856 119200 115528
rect 1025 114576 119120 114856
rect 1025 113904 119200 114576
rect 1025 113624 119120 113904
rect 1025 112952 119200 113624
rect 1025 112672 119120 112952
rect 1025 112000 119200 112672
rect 1025 111720 119120 112000
rect 1025 111184 119200 111720
rect 1025 110904 119120 111184
rect 1025 110232 119200 110904
rect 1025 109952 119120 110232
rect 1025 109280 119200 109952
rect 1025 109000 119120 109280
rect 1025 108328 119200 109000
rect 1025 108048 119120 108328
rect 1025 107376 119200 108048
rect 1025 107096 119120 107376
rect 1025 106424 119200 107096
rect 1025 106144 119120 106424
rect 1025 105472 119200 106144
rect 1025 105192 119120 105472
rect 1025 104520 119200 105192
rect 1025 104240 119120 104520
rect 1025 103568 119200 104240
rect 1025 103288 119120 103568
rect 1025 102752 119200 103288
rect 1025 102472 119120 102752
rect 1025 101800 119200 102472
rect 1025 101520 119120 101800
rect 1025 100848 119200 101520
rect 1025 100568 119120 100848
rect 1025 99896 119200 100568
rect 1025 99616 119120 99896
rect 1025 98944 119200 99616
rect 1025 98664 119120 98944
rect 1025 97992 119200 98664
rect 1025 97712 119120 97992
rect 1025 97040 119200 97712
rect 1025 96760 119120 97040
rect 1025 96088 119200 96760
rect 1025 95808 119120 96088
rect 1025 95136 119200 95808
rect 1025 94856 119120 95136
rect 1025 94320 119200 94856
rect 1025 94040 119120 94320
rect 1025 93368 119200 94040
rect 1025 93088 119120 93368
rect 1025 92416 119200 93088
rect 1025 92136 119120 92416
rect 1025 91464 119200 92136
rect 1025 91184 119120 91464
rect 1025 90512 119200 91184
rect 1025 90232 119120 90512
rect 1025 89560 119200 90232
rect 1025 89280 119120 89560
rect 1025 88608 119200 89280
rect 1025 88328 119120 88608
rect 1025 87656 119200 88328
rect 1025 87376 119120 87656
rect 1025 86704 119200 87376
rect 1025 86424 119120 86704
rect 1025 85888 119200 86424
rect 1025 85608 119120 85888
rect 1025 84936 119200 85608
rect 1025 84656 119120 84936
rect 1025 83984 119200 84656
rect 1025 83704 119120 83984
rect 1025 83032 119200 83704
rect 1025 82752 119120 83032
rect 1025 82080 119200 82752
rect 1025 81800 119120 82080
rect 1025 81128 119200 81800
rect 1025 80848 119120 81128
rect 1025 80176 119200 80848
rect 1025 79896 119120 80176
rect 1025 79224 119200 79896
rect 1025 78944 119120 79224
rect 1025 78272 119200 78944
rect 1025 77992 119120 78272
rect 1025 77456 119200 77992
rect 1025 77176 119120 77456
rect 1025 76504 119200 77176
rect 1025 76224 119120 76504
rect 1025 75552 119200 76224
rect 1025 75272 119120 75552
rect 1025 74600 119200 75272
rect 1025 74320 119120 74600
rect 1025 73648 119200 74320
rect 1025 73368 119120 73648
rect 1025 72696 119200 73368
rect 1025 72416 119120 72696
rect 1025 71744 119200 72416
rect 1025 71464 119120 71744
rect 1025 70792 119200 71464
rect 1025 70512 119120 70792
rect 1025 69840 119200 70512
rect 1025 69560 119120 69840
rect 1025 69024 119200 69560
rect 1025 68744 119120 69024
rect 1025 68072 119200 68744
rect 1025 67792 119120 68072
rect 1025 67120 119200 67792
rect 1025 66840 119120 67120
rect 1025 66168 119200 66840
rect 1025 65888 119120 66168
rect 1025 65216 119200 65888
rect 1025 64936 119120 65216
rect 1025 64264 119200 64936
rect 1025 63984 119120 64264
rect 1025 63312 119200 63984
rect 1025 63032 119120 63312
rect 1025 62360 119200 63032
rect 1025 62080 119120 62360
rect 1025 61408 119200 62080
rect 1025 61128 119120 61408
rect 1025 60592 119200 61128
rect 1025 60312 119120 60592
rect 1025 59640 119200 60312
rect 1025 59360 119120 59640
rect 1025 58688 119200 59360
rect 1025 58408 119120 58688
rect 1025 57736 119200 58408
rect 1025 57456 119120 57736
rect 1025 56784 119200 57456
rect 1025 56504 119120 56784
rect 1025 55832 119200 56504
rect 1025 55552 119120 55832
rect 1025 54880 119200 55552
rect 1025 54600 119120 54880
rect 1025 53928 119200 54600
rect 1025 53648 119120 53928
rect 1025 52976 119200 53648
rect 1025 52696 119120 52976
rect 1025 52024 119200 52696
rect 1025 51744 119120 52024
rect 1025 51208 119200 51744
rect 1025 50928 119120 51208
rect 1025 50256 119200 50928
rect 1025 49976 119120 50256
rect 1025 49304 119200 49976
rect 1025 49024 119120 49304
rect 1025 48352 119200 49024
rect 1025 48072 119120 48352
rect 1025 47400 119200 48072
rect 1025 47120 119120 47400
rect 1025 46448 119200 47120
rect 1025 46168 119120 46448
rect 1025 45496 119200 46168
rect 1025 45216 119120 45496
rect 1025 44544 119200 45216
rect 1025 44264 119120 44544
rect 1025 43592 119200 44264
rect 1025 43312 119120 43592
rect 1025 42776 119200 43312
rect 1025 42496 119120 42776
rect 1025 41824 119200 42496
rect 1025 41544 119120 41824
rect 1025 40872 119200 41544
rect 1025 40592 119120 40872
rect 1025 39920 119200 40592
rect 1025 39640 119120 39920
rect 1025 38968 119200 39640
rect 1025 38688 119120 38968
rect 1025 38016 119200 38688
rect 1025 37736 119120 38016
rect 1025 37064 119200 37736
rect 1025 36784 119120 37064
rect 1025 36112 119200 36784
rect 1025 35832 119120 36112
rect 1025 35160 119200 35832
rect 1025 34880 119120 35160
rect 1025 34344 119200 34880
rect 1025 34064 119120 34344
rect 1025 33392 119200 34064
rect 1025 33112 119120 33392
rect 1025 32440 119200 33112
rect 1025 32160 119120 32440
rect 1025 31488 119200 32160
rect 1025 31208 119120 31488
rect 1025 30536 119200 31208
rect 1025 30256 119120 30536
rect 1025 29584 119200 30256
rect 1025 29304 119120 29584
rect 1025 28632 119200 29304
rect 1025 28352 119120 28632
rect 1025 27680 119200 28352
rect 1025 27400 119120 27680
rect 1025 26728 119200 27400
rect 1025 26448 119120 26728
rect 1025 25912 119200 26448
rect 1025 25632 119120 25912
rect 1025 24960 119200 25632
rect 1025 24680 119120 24960
rect 1025 24008 119200 24680
rect 1025 23728 119120 24008
rect 1025 23056 119200 23728
rect 1025 22776 119120 23056
rect 1025 22104 119200 22776
rect 1025 21824 119120 22104
rect 1025 21152 119200 21824
rect 1025 20872 119120 21152
rect 1025 20200 119200 20872
rect 1025 19920 119120 20200
rect 1025 19248 119200 19920
rect 1025 18968 119120 19248
rect 1025 18296 119200 18968
rect 1025 18016 119120 18296
rect 1025 17480 119200 18016
rect 1025 17200 119120 17480
rect 1025 16528 119200 17200
rect 1025 16248 119120 16528
rect 1025 15576 119200 16248
rect 1025 15296 119120 15576
rect 1025 14624 119200 15296
rect 1025 14344 119120 14624
rect 1025 13672 119200 14344
rect 1025 13392 119120 13672
rect 1025 12720 119200 13392
rect 1025 12440 119120 12720
rect 1025 11768 119200 12440
rect 1025 11488 119120 11768
rect 1025 10816 119200 11488
rect 1025 10536 119120 10816
rect 1025 9864 119200 10536
rect 1025 9584 119120 9864
rect 1025 9048 119200 9584
rect 1025 8768 119120 9048
rect 1025 8096 119200 8768
rect 1025 7816 119120 8096
rect 1025 7144 119200 7816
rect 1025 6864 119120 7144
rect 1025 6192 119200 6864
rect 1025 5912 119120 6192
rect 1025 5240 119200 5912
rect 1025 4960 119120 5240
rect 1025 4288 119200 4960
rect 1025 4008 119120 4288
rect 1025 3336 119200 4008
rect 1025 3056 119120 3336
rect 1025 2384 119200 3056
rect 1025 2104 119120 2384
rect 1025 1432 119200 2104
rect 1025 1152 119120 1432
rect 1025 616 119200 1152
rect 1025 446 119120 616
<< metal4 >>
rect 1794 2128 2414 117552
rect 19794 2128 20414 117552
rect 37794 2128 38414 117552
rect 55794 2128 56414 117552
rect 73794 2128 74414 117552
rect 91794 2128 92414 117552
rect 109794 2128 110414 117552
<< obsm4 >>
rect 1531 2347 1714 113525
rect 2494 2347 19714 113525
rect 20494 2347 37714 113525
rect 38494 2347 55714 113525
rect 56494 2347 73714 113525
rect 74494 2347 91714 113525
rect 92494 2347 109714 113525
rect 110494 2347 116781 113525
<< labels >>
rlabel metal4 s 19794 2128 20414 117552 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 55794 2128 56414 117552 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 91794 2128 92414 117552 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1794 2128 2414 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 37794 2128 38414 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 73794 2128 74414 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 109794 2128 110414 117552 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 119200 416 120000 536 6 a[0]
port 3 nsew signal input
rlabel metal3 s 119200 9664 120000 9784 6 a[10]
port 4 nsew signal input
rlabel metal3 s 119200 10616 120000 10736 6 a[11]
port 5 nsew signal input
rlabel metal3 s 119200 11568 120000 11688 6 a[12]
port 6 nsew signal input
rlabel metal3 s 119200 12520 120000 12640 6 a[13]
port 7 nsew signal input
rlabel metal3 s 119200 13472 120000 13592 6 a[14]
port 8 nsew signal input
rlabel metal3 s 119200 14424 120000 14544 6 a[15]
port 9 nsew signal input
rlabel metal3 s 119200 15376 120000 15496 6 a[16]
port 10 nsew signal input
rlabel metal3 s 119200 16328 120000 16448 6 a[17]
port 11 nsew signal input
rlabel metal3 s 119200 17280 120000 17400 6 a[18]
port 12 nsew signal input
rlabel metal3 s 119200 18096 120000 18216 6 a[19]
port 13 nsew signal input
rlabel metal3 s 119200 1232 120000 1352 6 a[1]
port 14 nsew signal input
rlabel metal3 s 119200 19048 120000 19168 6 a[20]
port 15 nsew signal input
rlabel metal3 s 119200 20000 120000 20120 6 a[21]
port 16 nsew signal input
rlabel metal3 s 119200 20952 120000 21072 6 a[22]
port 17 nsew signal input
rlabel metal3 s 119200 21904 120000 22024 6 a[23]
port 18 nsew signal input
rlabel metal3 s 119200 22856 120000 22976 6 a[24]
port 19 nsew signal input
rlabel metal3 s 119200 23808 120000 23928 6 a[25]
port 20 nsew signal input
rlabel metal3 s 119200 24760 120000 24880 6 a[26]
port 21 nsew signal input
rlabel metal3 s 119200 25712 120000 25832 6 a[27]
port 22 nsew signal input
rlabel metal3 s 119200 26528 120000 26648 6 a[28]
port 23 nsew signal input
rlabel metal3 s 119200 27480 120000 27600 6 a[29]
port 24 nsew signal input
rlabel metal3 s 119200 2184 120000 2304 6 a[2]
port 25 nsew signal input
rlabel metal3 s 119200 28432 120000 28552 6 a[30]
port 26 nsew signal input
rlabel metal3 s 119200 29384 120000 29504 6 a[31]
port 27 nsew signal input
rlabel metal3 s 119200 30336 120000 30456 6 a[32]
port 28 nsew signal input
rlabel metal3 s 119200 31288 120000 31408 6 a[33]
port 29 nsew signal input
rlabel metal3 s 119200 32240 120000 32360 6 a[34]
port 30 nsew signal input
rlabel metal3 s 119200 33192 120000 33312 6 a[35]
port 31 nsew signal input
rlabel metal3 s 119200 34144 120000 34264 6 a[36]
port 32 nsew signal input
rlabel metal3 s 119200 34960 120000 35080 6 a[37]
port 33 nsew signal input
rlabel metal3 s 119200 35912 120000 36032 6 a[38]
port 34 nsew signal input
rlabel metal3 s 119200 36864 120000 36984 6 a[39]
port 35 nsew signal input
rlabel metal3 s 119200 3136 120000 3256 6 a[3]
port 36 nsew signal input
rlabel metal3 s 119200 37816 120000 37936 6 a[40]
port 37 nsew signal input
rlabel metal3 s 119200 38768 120000 38888 6 a[41]
port 38 nsew signal input
rlabel metal3 s 119200 39720 120000 39840 6 a[42]
port 39 nsew signal input
rlabel metal3 s 119200 40672 120000 40792 6 a[43]
port 40 nsew signal input
rlabel metal3 s 119200 41624 120000 41744 6 a[44]
port 41 nsew signal input
rlabel metal3 s 119200 42576 120000 42696 6 a[45]
port 42 nsew signal input
rlabel metal3 s 119200 43392 120000 43512 6 a[46]
port 43 nsew signal input
rlabel metal3 s 119200 44344 120000 44464 6 a[47]
port 44 nsew signal input
rlabel metal3 s 119200 45296 120000 45416 6 a[48]
port 45 nsew signal input
rlabel metal3 s 119200 46248 120000 46368 6 a[49]
port 46 nsew signal input
rlabel metal3 s 119200 4088 120000 4208 6 a[4]
port 47 nsew signal input
rlabel metal3 s 119200 47200 120000 47320 6 a[50]
port 48 nsew signal input
rlabel metal3 s 119200 48152 120000 48272 6 a[51]
port 49 nsew signal input
rlabel metal3 s 119200 49104 120000 49224 6 a[52]
port 50 nsew signal input
rlabel metal3 s 119200 50056 120000 50176 6 a[53]
port 51 nsew signal input
rlabel metal3 s 119200 51008 120000 51128 6 a[54]
port 52 nsew signal input
rlabel metal3 s 119200 51824 120000 51944 6 a[55]
port 53 nsew signal input
rlabel metal3 s 119200 52776 120000 52896 6 a[56]
port 54 nsew signal input
rlabel metal3 s 119200 53728 120000 53848 6 a[57]
port 55 nsew signal input
rlabel metal3 s 119200 54680 120000 54800 6 a[58]
port 56 nsew signal input
rlabel metal3 s 119200 55632 120000 55752 6 a[59]
port 57 nsew signal input
rlabel metal3 s 119200 5040 120000 5160 6 a[5]
port 58 nsew signal input
rlabel metal3 s 119200 56584 120000 56704 6 a[60]
port 59 nsew signal input
rlabel metal3 s 119200 57536 120000 57656 6 a[61]
port 60 nsew signal input
rlabel metal3 s 119200 58488 120000 58608 6 a[62]
port 61 nsew signal input
rlabel metal3 s 119200 59440 120000 59560 6 a[63]
port 62 nsew signal input
rlabel metal3 s 119200 5992 120000 6112 6 a[6]
port 63 nsew signal input
rlabel metal3 s 119200 6944 120000 7064 6 a[7]
port 64 nsew signal input
rlabel metal3 s 119200 7896 120000 8016 6 a[8]
port 65 nsew signal input
rlabel metal3 s 119200 8848 120000 8968 6 a[9]
port 66 nsew signal input
rlabel metal3 s 119200 60392 120000 60512 6 b[0]
port 67 nsew signal input
rlabel metal3 s 119200 69640 120000 69760 6 b[10]
port 68 nsew signal input
rlabel metal3 s 119200 70592 120000 70712 6 b[11]
port 69 nsew signal input
rlabel metal3 s 119200 71544 120000 71664 6 b[12]
port 70 nsew signal input
rlabel metal3 s 119200 72496 120000 72616 6 b[13]
port 71 nsew signal input
rlabel metal3 s 119200 73448 120000 73568 6 b[14]
port 72 nsew signal input
rlabel metal3 s 119200 74400 120000 74520 6 b[15]
port 73 nsew signal input
rlabel metal3 s 119200 75352 120000 75472 6 b[16]
port 74 nsew signal input
rlabel metal3 s 119200 76304 120000 76424 6 b[17]
port 75 nsew signal input
rlabel metal3 s 119200 77256 120000 77376 6 b[18]
port 76 nsew signal input
rlabel metal3 s 119200 78072 120000 78192 6 b[19]
port 77 nsew signal input
rlabel metal3 s 119200 61208 120000 61328 6 b[1]
port 78 nsew signal input
rlabel metal3 s 119200 79024 120000 79144 6 b[20]
port 79 nsew signal input
rlabel metal3 s 119200 79976 120000 80096 6 b[21]
port 80 nsew signal input
rlabel metal3 s 119200 80928 120000 81048 6 b[22]
port 81 nsew signal input
rlabel metal3 s 119200 81880 120000 82000 6 b[23]
port 82 nsew signal input
rlabel metal3 s 119200 82832 120000 82952 6 b[24]
port 83 nsew signal input
rlabel metal3 s 119200 83784 120000 83904 6 b[25]
port 84 nsew signal input
rlabel metal3 s 119200 84736 120000 84856 6 b[26]
port 85 nsew signal input
rlabel metal3 s 119200 85688 120000 85808 6 b[27]
port 86 nsew signal input
rlabel metal3 s 119200 86504 120000 86624 6 b[28]
port 87 nsew signal input
rlabel metal3 s 119200 87456 120000 87576 6 b[29]
port 88 nsew signal input
rlabel metal3 s 119200 62160 120000 62280 6 b[2]
port 89 nsew signal input
rlabel metal3 s 119200 88408 120000 88528 6 b[30]
port 90 nsew signal input
rlabel metal3 s 119200 89360 120000 89480 6 b[31]
port 91 nsew signal input
rlabel metal3 s 119200 90312 120000 90432 6 b[32]
port 92 nsew signal input
rlabel metal3 s 119200 91264 120000 91384 6 b[33]
port 93 nsew signal input
rlabel metal3 s 119200 92216 120000 92336 6 b[34]
port 94 nsew signal input
rlabel metal3 s 119200 93168 120000 93288 6 b[35]
port 95 nsew signal input
rlabel metal3 s 119200 94120 120000 94240 6 b[36]
port 96 nsew signal input
rlabel metal3 s 119200 94936 120000 95056 6 b[37]
port 97 nsew signal input
rlabel metal3 s 119200 95888 120000 96008 6 b[38]
port 98 nsew signal input
rlabel metal3 s 119200 96840 120000 96960 6 b[39]
port 99 nsew signal input
rlabel metal3 s 119200 63112 120000 63232 6 b[3]
port 100 nsew signal input
rlabel metal3 s 119200 97792 120000 97912 6 b[40]
port 101 nsew signal input
rlabel metal3 s 119200 98744 120000 98864 6 b[41]
port 102 nsew signal input
rlabel metal3 s 119200 99696 120000 99816 6 b[42]
port 103 nsew signal input
rlabel metal3 s 119200 100648 120000 100768 6 b[43]
port 104 nsew signal input
rlabel metal3 s 119200 101600 120000 101720 6 b[44]
port 105 nsew signal input
rlabel metal3 s 119200 102552 120000 102672 6 b[45]
port 106 nsew signal input
rlabel metal3 s 119200 103368 120000 103488 6 b[46]
port 107 nsew signal input
rlabel metal3 s 119200 104320 120000 104440 6 b[47]
port 108 nsew signal input
rlabel metal3 s 119200 105272 120000 105392 6 b[48]
port 109 nsew signal input
rlabel metal3 s 119200 106224 120000 106344 6 b[49]
port 110 nsew signal input
rlabel metal3 s 119200 64064 120000 64184 6 b[4]
port 111 nsew signal input
rlabel metal3 s 119200 107176 120000 107296 6 b[50]
port 112 nsew signal input
rlabel metal3 s 119200 108128 120000 108248 6 b[51]
port 113 nsew signal input
rlabel metal3 s 119200 109080 120000 109200 6 b[52]
port 114 nsew signal input
rlabel metal3 s 119200 110032 120000 110152 6 b[53]
port 115 nsew signal input
rlabel metal3 s 119200 110984 120000 111104 6 b[54]
port 116 nsew signal input
rlabel metal3 s 119200 111800 120000 111920 6 b[55]
port 117 nsew signal input
rlabel metal3 s 119200 112752 120000 112872 6 b[56]
port 118 nsew signal input
rlabel metal3 s 119200 113704 120000 113824 6 b[57]
port 119 nsew signal input
rlabel metal3 s 119200 114656 120000 114776 6 b[58]
port 120 nsew signal input
rlabel metal3 s 119200 115608 120000 115728 6 b[59]
port 121 nsew signal input
rlabel metal3 s 119200 65016 120000 65136 6 b[5]
port 122 nsew signal input
rlabel metal3 s 119200 116560 120000 116680 6 b[60]
port 123 nsew signal input
rlabel metal3 s 119200 117512 120000 117632 6 b[61]
port 124 nsew signal input
rlabel metal3 s 119200 118464 120000 118584 6 b[62]
port 125 nsew signal input
rlabel metal3 s 119200 119416 120000 119536 6 b[63]
port 126 nsew signal input
rlabel metal3 s 119200 65968 120000 66088 6 b[6]
port 127 nsew signal input
rlabel metal3 s 119200 66920 120000 67040 6 b[7]
port 128 nsew signal input
rlabel metal3 s 119200 67872 120000 67992 6 b[8]
port 129 nsew signal input
rlabel metal3 s 119200 68824 120000 68944 6 b[9]
port 130 nsew signal input
rlabel metal2 s 478 0 534 800 6 c[0]
port 131 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 c[100]
port 132 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 c[101]
port 133 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 c[102]
port 134 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 c[103]
port 135 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 c[104]
port 136 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 c[105]
port 137 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 c[106]
port 138 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 c[107]
port 139 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 c[108]
port 140 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 c[109]
port 141 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 c[10]
port 142 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 c[110]
port 143 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 c[111]
port 144 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 c[112]
port 145 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 c[113]
port 146 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 c[114]
port 147 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 c[115]
port 148 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 c[116]
port 149 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 c[117]
port 150 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 c[118]
port 151 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 c[119]
port 152 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 c[11]
port 153 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 c[120]
port 154 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 c[121]
port 155 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 c[122]
port 156 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 c[123]
port 157 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 c[124]
port 158 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 c[125]
port 159 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 c[126]
port 160 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 c[127]
port 161 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 c[12]
port 162 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 c[13]
port 163 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 c[14]
port 164 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 c[15]
port 165 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 c[16]
port 166 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 c[17]
port 167 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 c[18]
port 168 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 c[19]
port 169 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 c[1]
port 170 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 c[20]
port 171 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 c[21]
port 172 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 c[22]
port 173 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 c[23]
port 174 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 c[24]
port 175 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 c[25]
port 176 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 c[26]
port 177 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 c[27]
port 178 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 c[28]
port 179 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 c[29]
port 180 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 c[2]
port 181 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 c[30]
port 182 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 c[31]
port 183 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 c[32]
port 184 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 c[33]
port 185 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 c[34]
port 186 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 c[35]
port 187 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 c[36]
port 188 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 c[37]
port 189 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 c[38]
port 190 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 c[39]
port 191 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 c[3]
port 192 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 c[40]
port 193 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 c[41]
port 194 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 c[42]
port 195 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 c[43]
port 196 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 c[44]
port 197 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 c[45]
port 198 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 c[46]
port 199 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 c[47]
port 200 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 c[48]
port 201 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 c[49]
port 202 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 c[4]
port 203 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 c[50]
port 204 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 c[51]
port 205 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 c[52]
port 206 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 c[53]
port 207 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 c[54]
port 208 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 c[55]
port 209 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 c[56]
port 210 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 c[57]
port 211 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 c[58]
port 212 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 c[59]
port 213 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 c[5]
port 214 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 c[60]
port 215 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 c[61]
port 216 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 c[62]
port 217 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 c[63]
port 218 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 c[64]
port 219 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 c[65]
port 220 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 c[66]
port 221 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 c[67]
port 222 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 c[68]
port 223 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 c[69]
port 224 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 c[6]
port 225 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 c[70]
port 226 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 c[71]
port 227 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 c[72]
port 228 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 c[73]
port 229 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 c[74]
port 230 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 c[75]
port 231 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 c[76]
port 232 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 c[77]
port 233 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 c[78]
port 234 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 c[79]
port 235 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 c[7]
port 236 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 c[80]
port 237 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 c[81]
port 238 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 c[82]
port 239 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 c[83]
port 240 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 c[84]
port 241 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 c[85]
port 242 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 c[86]
port 243 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 c[87]
port 244 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 c[88]
port 245 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 c[89]
port 246 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 c[8]
port 247 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 c[90]
port 248 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 c[91]
port 249 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 c[92]
port 250 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 c[93]
port 251 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 c[94]
port 252 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 c[95]
port 253 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 c[96]
port 254 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 c[97]
port 255 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 c[98]
port 256 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 c[99]
port 257 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 c[9]
port 258 nsew signal input
rlabel metal2 s 119434 119200 119490 120000 6 clk
port 259 nsew signal input
rlabel metal2 s 478 119200 534 120000 6 o[0]
port 260 nsew signal output
rlabel metal2 s 92754 119200 92810 120000 6 o[100]
port 261 nsew signal output
rlabel metal2 s 93674 119200 93730 120000 6 o[101]
port 262 nsew signal output
rlabel metal2 s 94594 119200 94650 120000 6 o[102]
port 263 nsew signal output
rlabel metal2 s 95514 119200 95570 120000 6 o[103]
port 264 nsew signal output
rlabel metal2 s 96434 119200 96490 120000 6 o[104]
port 265 nsew signal output
rlabel metal2 s 97354 119200 97410 120000 6 o[105]
port 266 nsew signal output
rlabel metal2 s 98274 119200 98330 120000 6 o[106]
port 267 nsew signal output
rlabel metal2 s 99194 119200 99250 120000 6 o[107]
port 268 nsew signal output
rlabel metal2 s 100114 119200 100170 120000 6 o[108]
port 269 nsew signal output
rlabel metal2 s 101034 119200 101090 120000 6 o[109]
port 270 nsew signal output
rlabel metal2 s 9678 119200 9734 120000 6 o[10]
port 271 nsew signal output
rlabel metal2 s 101954 119200 102010 120000 6 o[110]
port 272 nsew signal output
rlabel metal2 s 102874 119200 102930 120000 6 o[111]
port 273 nsew signal output
rlabel metal2 s 103794 119200 103850 120000 6 o[112]
port 274 nsew signal output
rlabel metal2 s 104714 119200 104770 120000 6 o[113]
port 275 nsew signal output
rlabel metal2 s 105634 119200 105690 120000 6 o[114]
port 276 nsew signal output
rlabel metal2 s 106554 119200 106610 120000 6 o[115]
port 277 nsew signal output
rlabel metal2 s 107474 119200 107530 120000 6 o[116]
port 278 nsew signal output
rlabel metal2 s 108394 119200 108450 120000 6 o[117]
port 279 nsew signal output
rlabel metal2 s 109314 119200 109370 120000 6 o[118]
port 280 nsew signal output
rlabel metal2 s 110234 119200 110290 120000 6 o[119]
port 281 nsew signal output
rlabel metal2 s 10598 119200 10654 120000 6 o[11]
port 282 nsew signal output
rlabel metal2 s 111154 119200 111210 120000 6 o[120]
port 283 nsew signal output
rlabel metal2 s 112074 119200 112130 120000 6 o[121]
port 284 nsew signal output
rlabel metal2 s 112994 119200 113050 120000 6 o[122]
port 285 nsew signal output
rlabel metal2 s 113914 119200 113970 120000 6 o[123]
port 286 nsew signal output
rlabel metal2 s 114834 119200 114890 120000 6 o[124]
port 287 nsew signal output
rlabel metal2 s 115754 119200 115810 120000 6 o[125]
port 288 nsew signal output
rlabel metal2 s 116674 119200 116730 120000 6 o[126]
port 289 nsew signal output
rlabel metal2 s 117594 119200 117650 120000 6 o[127]
port 290 nsew signal output
rlabel metal2 s 11518 119200 11574 120000 6 o[12]
port 291 nsew signal output
rlabel metal2 s 12438 119200 12494 120000 6 o[13]
port 292 nsew signal output
rlabel metal2 s 13358 119200 13414 120000 6 o[14]
port 293 nsew signal output
rlabel metal2 s 14278 119200 14334 120000 6 o[15]
port 294 nsew signal output
rlabel metal2 s 15198 119200 15254 120000 6 o[16]
port 295 nsew signal output
rlabel metal2 s 16118 119200 16174 120000 6 o[17]
port 296 nsew signal output
rlabel metal2 s 17038 119200 17094 120000 6 o[18]
port 297 nsew signal output
rlabel metal2 s 17958 119200 18014 120000 6 o[19]
port 298 nsew signal output
rlabel metal2 s 1398 119200 1454 120000 6 o[1]
port 299 nsew signal output
rlabel metal2 s 18878 119200 18934 120000 6 o[20]
port 300 nsew signal output
rlabel metal2 s 19798 119200 19854 120000 6 o[21]
port 301 nsew signal output
rlabel metal2 s 20718 119200 20774 120000 6 o[22]
port 302 nsew signal output
rlabel metal2 s 21638 119200 21694 120000 6 o[23]
port 303 nsew signal output
rlabel metal2 s 22558 119200 22614 120000 6 o[24]
port 304 nsew signal output
rlabel metal2 s 23478 119200 23534 120000 6 o[25]
port 305 nsew signal output
rlabel metal2 s 24398 119200 24454 120000 6 o[26]
port 306 nsew signal output
rlabel metal2 s 25318 119200 25374 120000 6 o[27]
port 307 nsew signal output
rlabel metal2 s 26238 119200 26294 120000 6 o[28]
port 308 nsew signal output
rlabel metal2 s 27158 119200 27214 120000 6 o[29]
port 309 nsew signal output
rlabel metal2 s 2318 119200 2374 120000 6 o[2]
port 310 nsew signal output
rlabel metal2 s 28078 119200 28134 120000 6 o[30]
port 311 nsew signal output
rlabel metal2 s 28998 119200 29054 120000 6 o[31]
port 312 nsew signal output
rlabel metal2 s 29918 119200 29974 120000 6 o[32]
port 313 nsew signal output
rlabel metal2 s 30930 119200 30986 120000 6 o[33]
port 314 nsew signal output
rlabel metal2 s 31850 119200 31906 120000 6 o[34]
port 315 nsew signal output
rlabel metal2 s 32770 119200 32826 120000 6 o[35]
port 316 nsew signal output
rlabel metal2 s 33690 119200 33746 120000 6 o[36]
port 317 nsew signal output
rlabel metal2 s 34610 119200 34666 120000 6 o[37]
port 318 nsew signal output
rlabel metal2 s 35530 119200 35586 120000 6 o[38]
port 319 nsew signal output
rlabel metal2 s 36450 119200 36506 120000 6 o[39]
port 320 nsew signal output
rlabel metal2 s 3238 119200 3294 120000 6 o[3]
port 321 nsew signal output
rlabel metal2 s 37370 119200 37426 120000 6 o[40]
port 322 nsew signal output
rlabel metal2 s 38290 119200 38346 120000 6 o[41]
port 323 nsew signal output
rlabel metal2 s 39210 119200 39266 120000 6 o[42]
port 324 nsew signal output
rlabel metal2 s 40130 119200 40186 120000 6 o[43]
port 325 nsew signal output
rlabel metal2 s 41050 119200 41106 120000 6 o[44]
port 326 nsew signal output
rlabel metal2 s 41970 119200 42026 120000 6 o[45]
port 327 nsew signal output
rlabel metal2 s 42890 119200 42946 120000 6 o[46]
port 328 nsew signal output
rlabel metal2 s 43810 119200 43866 120000 6 o[47]
port 329 nsew signal output
rlabel metal2 s 44730 119200 44786 120000 6 o[48]
port 330 nsew signal output
rlabel metal2 s 45650 119200 45706 120000 6 o[49]
port 331 nsew signal output
rlabel metal2 s 4158 119200 4214 120000 6 o[4]
port 332 nsew signal output
rlabel metal2 s 46570 119200 46626 120000 6 o[50]
port 333 nsew signal output
rlabel metal2 s 47490 119200 47546 120000 6 o[51]
port 334 nsew signal output
rlabel metal2 s 48410 119200 48466 120000 6 o[52]
port 335 nsew signal output
rlabel metal2 s 49330 119200 49386 120000 6 o[53]
port 336 nsew signal output
rlabel metal2 s 50250 119200 50306 120000 6 o[54]
port 337 nsew signal output
rlabel metal2 s 51170 119200 51226 120000 6 o[55]
port 338 nsew signal output
rlabel metal2 s 52090 119200 52146 120000 6 o[56]
port 339 nsew signal output
rlabel metal2 s 53010 119200 53066 120000 6 o[57]
port 340 nsew signal output
rlabel metal2 s 53930 119200 53986 120000 6 o[58]
port 341 nsew signal output
rlabel metal2 s 54850 119200 54906 120000 6 o[59]
port 342 nsew signal output
rlabel metal2 s 5078 119200 5134 120000 6 o[5]
port 343 nsew signal output
rlabel metal2 s 55770 119200 55826 120000 6 o[60]
port 344 nsew signal output
rlabel metal2 s 56690 119200 56746 120000 6 o[61]
port 345 nsew signal output
rlabel metal2 s 57610 119200 57666 120000 6 o[62]
port 346 nsew signal output
rlabel metal2 s 58530 119200 58586 120000 6 o[63]
port 347 nsew signal output
rlabel metal2 s 59450 119200 59506 120000 6 o[64]
port 348 nsew signal output
rlabel metal2 s 60462 119200 60518 120000 6 o[65]
port 349 nsew signal output
rlabel metal2 s 61382 119200 61438 120000 6 o[66]
port 350 nsew signal output
rlabel metal2 s 62302 119200 62358 120000 6 o[67]
port 351 nsew signal output
rlabel metal2 s 63222 119200 63278 120000 6 o[68]
port 352 nsew signal output
rlabel metal2 s 64142 119200 64198 120000 6 o[69]
port 353 nsew signal output
rlabel metal2 s 5998 119200 6054 120000 6 o[6]
port 354 nsew signal output
rlabel metal2 s 65062 119200 65118 120000 6 o[70]
port 355 nsew signal output
rlabel metal2 s 65982 119200 66038 120000 6 o[71]
port 356 nsew signal output
rlabel metal2 s 66902 119200 66958 120000 6 o[72]
port 357 nsew signal output
rlabel metal2 s 67822 119200 67878 120000 6 o[73]
port 358 nsew signal output
rlabel metal2 s 68742 119200 68798 120000 6 o[74]
port 359 nsew signal output
rlabel metal2 s 69662 119200 69718 120000 6 o[75]
port 360 nsew signal output
rlabel metal2 s 70582 119200 70638 120000 6 o[76]
port 361 nsew signal output
rlabel metal2 s 71502 119200 71558 120000 6 o[77]
port 362 nsew signal output
rlabel metal2 s 72422 119200 72478 120000 6 o[78]
port 363 nsew signal output
rlabel metal2 s 73342 119200 73398 120000 6 o[79]
port 364 nsew signal output
rlabel metal2 s 6918 119200 6974 120000 6 o[7]
port 365 nsew signal output
rlabel metal2 s 74262 119200 74318 120000 6 o[80]
port 366 nsew signal output
rlabel metal2 s 75182 119200 75238 120000 6 o[81]
port 367 nsew signal output
rlabel metal2 s 76102 119200 76158 120000 6 o[82]
port 368 nsew signal output
rlabel metal2 s 77022 119200 77078 120000 6 o[83]
port 369 nsew signal output
rlabel metal2 s 77942 119200 77998 120000 6 o[84]
port 370 nsew signal output
rlabel metal2 s 78862 119200 78918 120000 6 o[85]
port 371 nsew signal output
rlabel metal2 s 79782 119200 79838 120000 6 o[86]
port 372 nsew signal output
rlabel metal2 s 80702 119200 80758 120000 6 o[87]
port 373 nsew signal output
rlabel metal2 s 81622 119200 81678 120000 6 o[88]
port 374 nsew signal output
rlabel metal2 s 82542 119200 82598 120000 6 o[89]
port 375 nsew signal output
rlabel metal2 s 7838 119200 7894 120000 6 o[8]
port 376 nsew signal output
rlabel metal2 s 83462 119200 83518 120000 6 o[90]
port 377 nsew signal output
rlabel metal2 s 84382 119200 84438 120000 6 o[91]
port 378 nsew signal output
rlabel metal2 s 85302 119200 85358 120000 6 o[92]
port 379 nsew signal output
rlabel metal2 s 86222 119200 86278 120000 6 o[93]
port 380 nsew signal output
rlabel metal2 s 87142 119200 87198 120000 6 o[94]
port 381 nsew signal output
rlabel metal2 s 88062 119200 88118 120000 6 o[95]
port 382 nsew signal output
rlabel metal2 s 88982 119200 89038 120000 6 o[96]
port 383 nsew signal output
rlabel metal2 s 89902 119200 89958 120000 6 o[97]
port 384 nsew signal output
rlabel metal2 s 90914 119200 90970 120000 6 o[98]
port 385 nsew signal output
rlabel metal2 s 91834 119200 91890 120000 6 o[99]
port 386 nsew signal output
rlabel metal2 s 8758 119200 8814 120000 6 o[9]
port 387 nsew signal output
rlabel metal2 s 118514 119200 118570 120000 6 rst
port 388 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35824944
string GDS_FILE /scratch/mpw6/caravel_user_project/openlane/multiply_add_64x64/runs/multiply_add_64x64/results/signoff/multiply_add_64x64.magic.gds
string GDS_START 289886
<< end >>

