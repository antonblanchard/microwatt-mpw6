* NGSPICE file created from multiply_add_64x64.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fa_1 abstract view
.subckt sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_1 abstract view
.subckt sky130_fd_sc_hd__ha_1 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fa_2 abstract view
.subckt sky130_fd_sc_hd__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ha_2 abstract view
.subckt sky130_fd_sc_hd__ha_2 A B VGND VNB VPB VPWR COUT SUM
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

.subckt multiply_add_64x64 VGND VPWR a[0] a[10] a[11] a[12] a[13] a[14] a[15] a[16]
+ a[17] a[18] a[19] a[1] a[20] a[21] a[22] a[23] a[24] a[25] a[26] a[27] a[28] a[29]
+ a[2] a[30] a[31] a[32] a[33] a[34] a[35] a[36] a[37] a[38] a[39] a[3] a[40] a[41]
+ a[42] a[43] a[44] a[45] a[46] a[47] a[48] a[49] a[4] a[50] a[51] a[52] a[53] a[54]
+ a[55] a[56] a[57] a[58] a[59] a[5] a[60] a[61] a[62] a[63] a[6] a[7] a[8] a[9] b[0]
+ b[10] b[11] b[12] b[13] b[14] b[15] b[16] b[17] b[18] b[19] b[1] b[20] b[21] b[22]
+ b[23] b[24] b[25] b[26] b[27] b[28] b[29] b[2] b[30] b[31] b[32] b[33] b[34] b[35]
+ b[36] b[37] b[38] b[39] b[3] b[40] b[41] b[42] b[43] b[44] b[45] b[46] b[47] b[48]
+ b[49] b[4] b[50] b[51] b[52] b[53] b[54] b[55] b[56] b[57] b[58] b[59] b[5] b[60]
+ b[61] b[62] b[63] b[6] b[7] b[8] b[9] c[0] c[100] c[101] c[102] c[103] c[104] c[105]
+ c[106] c[107] c[108] c[109] c[10] c[110] c[111] c[112] c[113] c[114] c[115] c[116]
+ c[117] c[118] c[119] c[11] c[120] c[121] c[122] c[123] c[124] c[125] c[126] c[127]
+ c[12] c[13] c[14] c[15] c[16] c[17] c[18] c[19] c[1] c[20] c[21] c[22] c[23] c[24]
+ c[25] c[26] c[27] c[28] c[29] c[2] c[30] c[31] c[32] c[33] c[34] c[35] c[36] c[37]
+ c[38] c[39] c[3] c[40] c[41] c[42] c[43] c[44] c[45] c[46] c[47] c[48] c[49] c[4]
+ c[50] c[51] c[52] c[53] c[54] c[55] c[56] c[57] c[58] c[59] c[5] c[60] c[61] c[62]
+ c[63] c[64] c[65] c[66] c[67] c[68] c[69] c[6] c[70] c[71] c[72] c[73] c[74] c[75]
+ c[76] c[77] c[78] c[79] c[7] c[80] c[81] c[82] c[83] c[84] c[85] c[86] c[87] c[88]
+ c[89] c[8] c[90] c[91] c[92] c[93] c[94] c[95] c[96] c[97] c[98] c[99] c[9] clk
+ o[0] o[100] o[101] o[102] o[103] o[104] o[105] o[106] o[107] o[108] o[109] o[10]
+ o[110] o[111] o[112] o[113] o[114] o[115] o[116] o[117] o[118] o[119] o[11] o[120]
+ o[121] o[122] o[123] o[124] o[125] o[126] o[127] o[12] o[13] o[14] o[15] o[16] o[17]
+ o[18] o[19] o[1] o[20] o[21] o[22] o[23] o[24] o[25] o[26] o[27] o[28] o[29] o[2]
+ o[30] o[31] o[32] o[33] o[34] o[35] o[36] o[37] o[38] o[39] o[3] o[40] o[41] o[42]
+ o[43] o[44] o[45] o[46] o[47] o[48] o[49] o[4] o[50] o[51] o[52] o[53] o[54] o[55]
+ o[56] o[57] o[58] o[59] o[5] o[60] o[61] o[62] o[63] o[64] o[65] o[66] o[67] o[68]
+ o[69] o[6] o[70] o[71] o[72] o[73] o[74] o[75] o[76] o[77] o[78] o[79] o[7] o[80]
+ o[81] o[82] o[83] o[84] o[85] o[86] o[87] o[88] o[89] o[8] o[90] o[91] o[92] o[93]
+ o[94] o[95] o[96] o[97] o[98] o[99] o[9] rst
Xdadda_fa_1_57_8 dadda_fa_1_57_8/A dadda_fa_1_57_8/B dadda_fa_1_57_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_58_3/A dadda_fa_3_57_0/A sky130_fd_sc_hd__fa_1
XFILLER_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_104_0 dadda_fa_2_104_0/A U$$2875/X U$$3008/X VGND VGND VPWR VPWR dadda_fa_3_105_2/CIN
+ dadda_fa_3_104_3/B sky130_fd_sc_hd__fa_1
XFILLER_211_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1290 U$$1290/A U$$1330/B VGND VGND VPWR VPWR U$$1290/X sky130_fd_sc_hd__xor2_1
XFILLER_206_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_90_2 U$$2581/X U$$2714/X U$$2847/X VGND VGND VPWR VPWR dadda_fa_2_91_4/CIN
+ dadda_fa_2_90_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_11_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_83_1 U$$1769/X U$$1902/X U$$2035/X VGND VGND VPWR VPWR dadda_fa_2_84_2/A
+ dadda_fa_2_83_4/B sky130_fd_sc_hd__fa_1
XFILLER_81_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_60_0 dadda_fa_4_60_0/A dadda_fa_4_60_0/B dadda_fa_4_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/A dadda_fa_5_60_1/A sky130_fd_sc_hd__fa_1
XFILLER_77_306 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_76_0 U$$1489/X U$$1622/X U$$1755/X VGND VGND VPWR VPWR dadda_fa_2_77_0/B
+ dadda_fa_2_76_3/B sky130_fd_sc_hd__fa_1
XFILLER_104_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_840 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3609 U$$3609/A U$$3609/B VGND VGND VPWR VPWR U$$3609/X sky130_fd_sc_hd__xor2_1
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2908 U$$2908/A U$$2996/B VGND VGND VPWR VPWR U$$2908/X sky130_fd_sc_hd__xor2_1
XFILLER_172_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_202 _199_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2919 U$$4289/A1 U$$2919/A2 U$$3058/A1 U$$2919/B2 VGND VGND VPWR VPWR U$$2920/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 _209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_224 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_5_124_1 U$$4511/X input156/X VGND VGND VPWR VPWR dadda_fa_6_125_0/CIN dadda_fa_7_124_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 _292_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 input128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_198_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 U$$2828/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_954 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_363_ _363_/CLK _363_/D VGND VGND VPWR VPWR _363_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_294_ _423_/CLK _294_/D VGND VGND VPWR VPWR _294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_98_1 dadda_fa_3_98_1/A dadda_fa_3_98_1/B dadda_fa_3_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_0/CIN dadda_fa_4_98_2/A sky130_fd_sc_hd__fa_1
XFILLER_115_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_75_0 dadda_fa_6_75_0/A dadda_fa_6_75_0/B dadda_fa_6_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_76_0/B dadda_fa_7_75_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$370 U$$916/B1 U$$378/A2 U$$920/A1 U$$378/B2 VGND VGND VPWR VPWR U$$371/A sky130_fd_sc_hd__a22o_1
XU$$381 U$$381/A U$$395/B VGND VGND VPWR VPWR U$$381/X sky130_fd_sc_hd__xor2_1
XFILLER_33_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$392 U$$392/A1 U$$394/A2 U$$942/A1 U$$394/B2 VGND VGND VPWR VPWR U$$393/A sky130_fd_sc_hd__a22o_1
XFILLER_44_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_93_0 U$$2853/X U$$2986/X U$$3119/X VGND VGND VPWR VPWR dadda_fa_3_94_0/B
+ dadda_fa_3_93_2/B sky130_fd_sc_hd__fa_1
XFILLER_173_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1270 U$$3836/A VGND VGND VPWR VPWR U$$3774/B sky130_fd_sc_hd__buf_6
Xrepeater1281 U$$945/B VGND VGND VPWR VPWR U$$951/B sky130_fd_sc_hd__buf_6
Xrepeater1292 U$$3643/B VGND VGND VPWR VPWR U$$3637/B sky130_fd_sc_hd__buf_6
XFILLER_102_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_6 dadda_fa_1_62_6/A dadda_fa_1_62_6/B dadda_fa_1_62_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_2/B dadda_fa_2_62_5/B sky130_fd_sc_hd__fa_1
XFILLER_68_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_55_5 U$$2777/X U$$2910/X U$$3043/X VGND VGND VPWR VPWR dadda_fa_2_56_2/A
+ dadda_fa_2_55_5/A sky130_fd_sc_hd__fa_1
XFILLER_67_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_48_4 U$$1699/X U$$1832/X U$$1965/X VGND VGND VPWR VPWR dadda_fa_2_49_2/B
+ dadda_fa_2_48_5/A sky130_fd_sc_hd__fa_1
XFILLER_83_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_18_2 dadda_fa_4_18_2/A dadda_fa_4_18_2/B dadda_ha_3_18_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_19_0/CIN dadda_fa_5_18_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_70_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_92_0 dadda_fa_7_92_0/A dadda_fa_7_92_0/B dadda_fa_7_92_0/CIN VGND VGND
+ VPWR VPWR _389_/D _260_/D sky130_fd_sc_hd__fa_1
XFILLER_17_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4107 U$$4242/B1 U$$4107/A2 U$$4107/B1 U$$4107/B2 VGND VGND VPWR VPWR U$$4108/A
+ sky130_fd_sc_hd__a22o_1
XU$$4118 U$$4392/A1 U$$4144/A2 U$$4394/A1 U$$4144/B2 VGND VGND VPWR VPWR U$$4119/A
+ sky130_fd_sc_hd__a22o_1
XU$$4129 U$$4129/A U$$4246/A VGND VGND VPWR VPWR U$$4129/X sky130_fd_sc_hd__xor2_1
XFILLER_77_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3406 U$$3817/A1 U$$3422/A2 U$$3545/A1 U$$3422/B2 VGND VGND VPWR VPWR U$$3407/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3417 U$$3417/A U$$3417/B VGND VGND VPWR VPWR U$$3417/X sky130_fd_sc_hd__xor2_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3428 U$$3510/B U$$3428/B VGND VGND VPWR VPWR U$$3428/X sky130_fd_sc_hd__and2_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3439 U$$3713/A1 U$$3527/A2 U$$3578/A1 U$$3527/B2 VGND VGND VPWR VPWR U$$3440/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2705 U$$2842/A1 U$$2607/X U$$2842/B1 U$$2608/X VGND VGND VPWR VPWR U$$2706/A sky130_fd_sc_hd__a22o_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2716 U$$2716/A U$$2716/B VGND VGND VPWR VPWR U$$2716/X sky130_fd_sc_hd__xor2_1
XFILLER_160_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2727 U$$3547/B1 U$$2727/A2 U$$3414/A1 U$$2727/B2 VGND VGND VPWR VPWR U$$2728/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2738 U$$2738/A U$$2739/A VGND VGND VPWR VPWR U$$2738/X sky130_fd_sc_hd__xor2_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2749 U$$2749/A U$$2755/B VGND VGND VPWR VPWR U$$2749/X sky130_fd_sc_hd__xor2_1
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_2 U$$845/X U$$978/X U$$1111/X VGND VGND VPWR VPWR dadda_fa_4_21_1/A
+ dadda_fa_4_20_2/B sky130_fd_sc_hd__fa_1
XFILLER_15_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_415_ _417_/CLK _415_/D VGND VGND VPWR VPWR _415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1023 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_346_ _351_/CLK _346_/D VGND VGND VPWR VPWR _346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1067 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_277_ _407_/CLK _277_/D VGND VGND VPWR VPWR _277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_72_5 dadda_fa_2_72_5/A dadda_fa_2_72_5/B dadda_fa_2_72_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_2/A dadda_fa_4_72_0/A sky130_fd_sc_hd__fa_1
XFILLER_190_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_65_4 dadda_fa_2_65_4/A dadda_fa_2_65_4/B dadda_fa_2_65_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/CIN dadda_fa_3_65_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_116_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater904 U$$4333/B1 VGND VGND VPWR VPWR U$$3922/B1 sky130_fd_sc_hd__buf_8
Xrepeater915 U$$3300/B1 VGND VGND VPWR VPWR U$$2343/A1 sky130_fd_sc_hd__buf_4
Xrepeater926 input97/X VGND VGND VPWR VPWR U$$4468/B1 sky130_fd_sc_hd__buf_4
XFILLER_56_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater937 input95/X VGND VGND VPWR VPWR U$$4055/A1 sky130_fd_sc_hd__buf_4
XFILLER_49_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_58_3 dadda_fa_2_58_3/A dadda_fa_2_58_3/B dadda_fa_2_58_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/B dadda_fa_3_58_3/B sky130_fd_sc_hd__fa_1
Xrepeater948 U$$4464/A1 VGND VGND VPWR VPWR U$$2957/A1 sky130_fd_sc_hd__buf_6
XFILLER_37_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater959 U$$2951/B1 VGND VGND VPWR VPWR U$$76/A1 sky130_fd_sc_hd__buf_6
XFILLER_37_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3940 U$$4488/A1 U$$3966/A2 U$$4077/B1 U$$3966/B2 VGND VGND VPWR VPWR U$$3941/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_28_1 dadda_fa_5_28_1/A dadda_fa_5_28_1/B dadda_fa_5_28_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_29_0/B dadda_fa_7_28_0/A sky130_fd_sc_hd__fa_2
XU$$3951 U$$3951/A U$$3972/A VGND VGND VPWR VPWR U$$3951/X sky130_fd_sc_hd__xor2_1
XFILLER_80_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3962 U$$4236/A1 U$$3966/A2 U$$4099/B1 U$$3966/B2 VGND VGND VPWR VPWR U$$3963/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3973 input53/X VGND VGND VPWR VPWR U$$3973/Y sky130_fd_sc_hd__inv_1
XU$$3984 U$$3984/A U$$4012/B VGND VGND VPWR VPWR U$$3984/X sky130_fd_sc_hd__xor2_1
XU$$3995 U$$4406/A1 U$$4035/A2 U$$4408/A1 U$$4035/B2 VGND VGND VPWR VPWR U$$3996/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_102_1 dadda_fa_5_102_1/A dadda_fa_5_102_1/B dadda_fa_5_102_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_103_0/B dadda_fa_7_102_0/A sky130_fd_sc_hd__fa_1
XFILLER_47_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput264 output264/A VGND VGND VPWR VPWR o[106] sky130_fd_sc_hd__buf_2
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput275 output275/A VGND VGND VPWR VPWR o[116] sky130_fd_sc_hd__buf_2
XFILLER_134_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput286 output286/A VGND VGND VPWR VPWR o[126] sky130_fd_sc_hd__buf_2
XFILLER_142_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput297 output297/A VGND VGND VPWR VPWR o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_60_3 U$$3186/X U$$3319/X U$$3452/X VGND VGND VPWR VPWR dadda_fa_2_61_1/B
+ dadda_fa_2_60_4/B sky130_fd_sc_hd__fa_1
XFILLER_114_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_53_2 U$$1177/X U$$1310/X U$$1443/X VGND VGND VPWR VPWR dadda_fa_2_54_1/A
+ dadda_fa_2_53_4/A sky130_fd_sc_hd__fa_1
XFILLER_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_30_1 dadda_fa_4_30_1/A dadda_fa_4_30_1/B dadda_fa_4_30_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/B dadda_fa_5_30_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_46_1 U$$498/X U$$631/X U$$764/X VGND VGND VPWR VPWR dadda_fa_2_47_2/A
+ dadda_fa_2_46_4/B sky130_fd_sc_hd__fa_2
XFILLER_167_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1034 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_23_0 dadda_fa_4_23_0/A dadda_fa_4_23_0/B dadda_fa_4_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/A dadda_fa_5_23_1/A sky130_fd_sc_hd__fa_1
XFILLER_71_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_39_0 U$$85/X U$$218/X U$$351/X VGND VGND VPWR VPWR dadda_fa_2_40_4/A dadda_fa_2_39_5/B
+ sky130_fd_sc_hd__fa_1
XFILLER_70_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_200_ _329_/CLK _200_/D VGND VGND VPWR VPWR _200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1105 final_adder.U$$174/B final_adder.U$$945/X VGND VGND VPWR VPWR
+ output364/A sky130_fd_sc_hd__xor2_1
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1116 final_adder.U$$162/A final_adder.U$$871/X VGND VGND VPWR VPWR
+ output376/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1127 final_adder.U$$152/B final_adder.U$$923/X VGND VGND VPWR VPWR
+ output261/A sky130_fd_sc_hd__xor2_2
XFILLER_7_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1138 final_adder.U$$140/A final_adder.U$$849/X VGND VGND VPWR VPWR
+ output273/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1149 final_adder.U$$130/B final_adder.U$$901/X VGND VGND VPWR VPWR
+ output285/A sky130_fd_sc_hd__xor2_1
XFILLER_164_450 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_75_3 dadda_fa_3_75_3/A dadda_fa_3_75_3/B dadda_fa_3_75_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_1/B dadda_fa_4_75_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_68_2 dadda_fa_3_68_2/A dadda_fa_3_68_2/B dadda_fa_3_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_1/A dadda_fa_4_68_2/B sky130_fd_sc_hd__fa_1
XFILLER_78_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_38_0 dadda_fa_6_38_0/A dadda_fa_6_38_0/B dadda_fa_6_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_39_0/B dadda_fa_7_38_0/CIN sky130_fd_sc_hd__fa_1
XU$$3203 U$$4297/B1 U$$3241/A2 U$$4162/B1 U$$3241/B2 VGND VGND VPWR VPWR U$$3204/A
+ sky130_fd_sc_hd__a22o_1
XU$$3214 U$$3214/A U$$3228/B VGND VGND VPWR VPWR U$$3214/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3225 U$$3908/B1 U$$3155/X input92/X U$$3156/X VGND VGND VPWR VPWR U$$3226/A sky130_fd_sc_hd__a22o_1
XFILLER_185_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3236 U$$3236/A U$$3242/B VGND VGND VPWR VPWR U$$3236/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$18 _314_/Q _186_/Q VGND VGND VPWR VPWR final_adder.U$$237/A2 final_adder.U$$236/A
+ sky130_fd_sc_hd__ha_1
XU$$3247 input103/X U$$3255/A2 U$$4480/B1 U$$3255/B2 VGND VGND VPWR VPWR U$$3248/A
+ sky130_fd_sc_hd__a22o_1
XU$$2502 U$$719/B1 U$$2596/A2 U$$312/A1 U$$2596/B2 VGND VGND VPWR VPWR U$$2503/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$29 _325_/Q _197_/Q VGND VGND VPWR VPWR final_adder.U$$227/B1 final_adder.U$$226/B
+ sky130_fd_sc_hd__ha_1
XU$$3258 U$$3258/A U$$3264/B VGND VGND VPWR VPWR U$$3258/X sky130_fd_sc_hd__xor2_1
XU$$2513 U$$2513/A U$$2597/B VGND VGND VPWR VPWR U$$2513/X sky130_fd_sc_hd__xor2_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2524 U$$3207/B1 U$$2524/A2 U$$2661/B1 U$$2524/B2 VGND VGND VPWR VPWR U$$2525/A
+ sky130_fd_sc_hd__a22o_1
XU$$3269 U$$3817/A1 U$$3277/A2 input116/X U$$3277/B2 VGND VGND VPWR VPWR U$$3270/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2535 U$$2535/A U$$2577/B VGND VGND VPWR VPWR U$$2535/X sky130_fd_sc_hd__xor2_1
XU$$2546 U$$2957/A1 U$$2558/A2 U$$3368/B1 U$$2558/B2 VGND VGND VPWR VPWR U$$2547/A
+ sky130_fd_sc_hd__a22o_1
XU$$1801 U$$979/A1 U$$1839/A2 U$$981/A1 U$$1839/B2 VGND VGND VPWR VPWR U$$1802/A sky130_fd_sc_hd__a22o_1
XU$$2557 U$$2557/A U$$2602/A VGND VGND VPWR VPWR U$$2557/X sky130_fd_sc_hd__xor2_1
XFILLER_34_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1812 U$$1812/A U$$1832/B VGND VGND VPWR VPWR U$$1812/X sky130_fd_sc_hd__xor2_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1823 U$$727/A1 U$$1869/A2 U$$727/B1 U$$1869/B2 VGND VGND VPWR VPWR U$$1824/A sky130_fd_sc_hd__a22o_1
XU$$2568 U$$2842/A1 U$$2470/X U$$2568/B1 U$$2471/X VGND VGND VPWR VPWR U$$2569/A sky130_fd_sc_hd__a22o_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2579 U$$2579/A U$$2603/A VGND VGND VPWR VPWR U$$2579/X sky130_fd_sc_hd__xor2_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1834 U$$1834/A U$$1840/B VGND VGND VPWR VPWR U$$1834/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1845 U$$3215/A1 U$$1879/A2 U$$1984/A1 U$$1879/B2 VGND VGND VPWR VPWR U$$1846/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1856 U$$1856/A U$$1880/B VGND VGND VPWR VPWR U$$1856/X sky130_fd_sc_hd__xor2_1
XU$$1867 U$$3235/B1 U$$1869/A2 U$$3376/A1 U$$1869/B2 VGND VGND VPWR VPWR U$$1868/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1878 U$$1878/A U$$1878/B VGND VGND VPWR VPWR U$$1878/X sky130_fd_sc_hd__xor2_1
XFILLER_202_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1889 U$$930/A1 U$$1915/A2 U$$2165/A1 U$$1915/B2 VGND VGND VPWR VPWR U$$1890/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_329_ _329_/CLK _329_/D VGND VGND VPWR VPWR _329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_3_1_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_192_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_70_2 dadda_fa_2_70_2/A dadda_fa_2_70_2/B dadda_fa_2_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/A dadda_fa_3_70_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_63_1 dadda_fa_2_63_1/A dadda_fa_2_63_1/B dadda_fa_2_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_0/CIN dadda_fa_3_63_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater701 U$$3978/X VGND VGND VPWR VPWR U$$4107/B2 sky130_fd_sc_hd__buf_6
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$508 final_adder.U$$516/B final_adder.U$$508/B VGND VGND VPWR VPWR
+ final_adder.U$$628/B sky130_fd_sc_hd__and2_1
Xrepeater712 U$$3819/B2 VGND VGND VPWR VPWR U$$3813/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$519 final_adder.U$$518/B final_adder.U$$403/X final_adder.U$$395/X
+ VGND VGND VPWR VPWR final_adder.U$$519/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_40_0 dadda_fa_5_40_0/A dadda_fa_5_40_0/B dadda_fa_5_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_41_0/A dadda_fa_6_40_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater723 U$$3644/B2 VGND VGND VPWR VPWR U$$3696/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_56_0 dadda_fa_2_56_0/A dadda_fa_2_56_0/B dadda_fa_2_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_0/B dadda_fa_3_56_2/B sky130_fd_sc_hd__fa_1
Xrepeater734 U$$3320/B2 VGND VGND VPWR VPWR U$$3394/B2 sky130_fd_sc_hd__buf_8
Xrepeater745 U$$3156/X VGND VGND VPWR VPWR U$$3227/B2 sky130_fd_sc_hd__buf_6
XFILLER_38_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater756 U$$3118/B2 VGND VGND VPWR VPWR U$$3082/B2 sky130_fd_sc_hd__buf_12
Xrepeater767 U$$340/B2 VGND VGND VPWR VPWR U$$316/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater778 U$$2858/B2 VGND VGND VPWR VPWR U$$2868/B2 sky130_fd_sc_hd__buf_4
XFILLER_49_191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4460 U$$4460/A1 U$$4388/X input93/X U$$4476/B2 VGND VGND VPWR VPWR U$$4461/A sky130_fd_sc_hd__a22o_1
XFILLER_93_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4471 U$$4471/A U$$4471/B VGND VGND VPWR VPWR U$$4471/X sky130_fd_sc_hd__xor2_1
Xrepeater789 U$$2711/B2 VGND VGND VPWR VPWR U$$2737/B2 sky130_fd_sc_hd__clkbuf_8
XU$$4482 input104/X U$$4388/X input105/X U$$4486/B2 VGND VGND VPWR VPWR U$$4483/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4493 U$$4493/A U$$4493/B VGND VGND VPWR VPWR U$$4493/X sky130_fd_sc_hd__xor2_1
XU$$3770 U$$3770/A U$$3774/B VGND VGND VPWR VPWR U$$3770/X sky130_fd_sc_hd__xor2_1
XU$$3781 input95/X U$$3819/A2 input96/X U$$3819/B2 VGND VGND VPWR VPWR U$$3782/A sky130_fd_sc_hd__a22o_1
XFILLER_64_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3792 U$$3792/A U$$3794/B VGND VGND VPWR VPWR U$$3792/X sky130_fd_sc_hd__xor2_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_450 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_85_2 dadda_fa_4_85_2/A dadda_fa_4_85_2/B dadda_fa_4_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/CIN dadda_fa_5_85_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_78_1 dadda_fa_4_78_1/A dadda_fa_4_78_1/B dadda_fa_4_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/B dadda_fa_5_78_1/B sky130_fd_sc_hd__fa_1
XFILLER_192_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_55_0 dadda_fa_7_55_0/A dadda_fa_7_55_0/B dadda_fa_7_55_0/CIN VGND VGND
+ VPWR VPWR _352_/D _223_/D sky130_fd_sc_hd__fa_1
XFILLER_115_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$903 U$$903/A U$$951/B VGND VGND VPWR VPWR U$$903/X sky130_fd_sc_hd__xor2_1
XU$$914 U$$914/A1 U$$918/A2 U$$914/B1 U$$918/B2 VGND VGND VPWR VPWR U$$915/A sky130_fd_sc_hd__a22o_1
XFILLER_44_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$925 U$$925/A U$$951/B VGND VGND VPWR VPWR U$$925/X sky130_fd_sc_hd__xor2_1
XU$$936 U$$936/A1 U$$826/X U$$936/B1 U$$827/X VGND VGND VPWR VPWR U$$937/A sky130_fd_sc_hd__a22o_1
XFILLER_71_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$947 U$$947/A U$$958/A VGND VGND VPWR VPWR U$$947/X sky130_fd_sc_hd__xor2_1
XFILLER_28_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$958 U$$958/A VGND VGND VPWR VPWR U$$958/Y sky130_fd_sc_hd__inv_1
XU$$969 U$$969/A1 U$$979/A2 U$$969/B1 U$$979/B2 VGND VGND VPWR VPWR U$$970/A sky130_fd_sc_hd__a22o_1
XU$$1108 U$$969/B1 U$$1138/A2 U$$2069/A1 U$$1138/B2 VGND VGND VPWR VPWR U$$1109/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1119 U$$1119/A U$$1137/B VGND VGND VPWR VPWR U$$1119/X sky130_fd_sc_hd__xor2_1
XFILLER_203_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_80_1 dadda_fa_3_80_1/A dadda_fa_3_80_1/B dadda_fa_3_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_0/CIN dadda_fa_4_80_2/A sky130_fd_sc_hd__fa_1
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_73_0 dadda_fa_3_73_0/A dadda_fa_3_73_0/B dadda_fa_3_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_0/B dadda_fa_4_73_1/CIN sky130_fd_sc_hd__fa_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3000 U$$3000/A U$$3013/A VGND VGND VPWR VPWR U$$3000/X sky130_fd_sc_hd__xor2_1
XU$$3011 U$$3557/B1 U$$3011/A2 U$$3011/B1 U$$3011/B2 VGND VGND VPWR VPWR U$$3012/A
+ sky130_fd_sc_hd__a22o_1
XU$$3022 U$$3159/A1 U$$3060/A2 U$$3159/B1 U$$3060/B2 VGND VGND VPWR VPWR U$$3023/A
+ sky130_fd_sc_hd__a22o_1
XU$$3033 U$$3033/A U$$3083/B VGND VGND VPWR VPWR U$$3033/X sky130_fd_sc_hd__xor2_1
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3044 U$$30/A1 U$$3124/A2 U$$32/A1 U$$3124/B2 VGND VGND VPWR VPWR U$$3045/A sky130_fd_sc_hd__a22o_1
XFILLER_47_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2310 U$$2445/B1 U$$2196/X U$$2312/A1 U$$2197/X VGND VGND VPWR VPWR U$$2311/A sky130_fd_sc_hd__a22o_1
XU$$3055 U$$3055/A U$$3075/B VGND VGND VPWR VPWR U$$3055/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_102_0 dadda_fa_4_102_0/A dadda_fa_4_102_0/B dadda_fa_4_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/A dadda_fa_5_102_1/A sky130_fd_sc_hd__fa_1
XU$$2321 U$$2321/A U$$2328/A VGND VGND VPWR VPWR U$$2321/X sky130_fd_sc_hd__xor2_1
XU$$3066 U$$4436/A1 U$$3108/A2 U$$4438/A1 U$$3108/B2 VGND VGND VPWR VPWR U$$3067/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_35_5 U$$2338/X input185/X dadda_fa_2_35_5/CIN VGND VGND VPWR VPWR dadda_fa_3_36_2/A
+ dadda_fa_4_35_0/A sky130_fd_sc_hd__fa_1
XU$$2332 input29/X U$$2332/B VGND VGND VPWR VPWR U$$2332/X sky130_fd_sc_hd__and2_1
XFILLER_62_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3077 U$$3077/A U$$3077/B VGND VGND VPWR VPWR U$$3077/X sky130_fd_sc_hd__xor2_1
XFILLER_35_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2343 U$$2343/A1 U$$2359/A2 U$$3987/B1 U$$2359/B2 VGND VGND VPWR VPWR U$$2344/A
+ sky130_fd_sc_hd__a22o_1
XU$$3088 U$$3088/A1 U$$3118/A2 U$$3499/B1 U$$3118/B2 VGND VGND VPWR VPWR U$$3089/A
+ sky130_fd_sc_hd__a22o_1
XU$$2354 U$$2354/A U$$2360/B VGND VGND VPWR VPWR U$$2354/X sky130_fd_sc_hd__xor2_1
XU$$3099 U$$3099/A U$$3109/B VGND VGND VPWR VPWR U$$3099/X sky130_fd_sc_hd__xor2_1
XFILLER_61_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1620 U$$1620/A U$$1620/B VGND VGND VPWR VPWR U$$1620/X sky130_fd_sc_hd__xor2_1
XFILLER_61_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2365 U$$995/A1 U$$2417/A2 U$$721/B1 U$$2417/B2 VGND VGND VPWR VPWR U$$2366/A sky130_fd_sc_hd__a22o_1
XU$$2376 U$$2376/A U$$2380/B VGND VGND VPWR VPWR U$$2376/X sky130_fd_sc_hd__xor2_1
XU$$1631 U$$2316/A1 U$$1637/A2 U$$4510/A1 U$$1637/B2 VGND VGND VPWR VPWR U$$1632/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1642 U$$1642/A U$$1644/A VGND VGND VPWR VPWR U$$1642/X sky130_fd_sc_hd__xor2_1
XU$$2387 U$$3207/B1 U$$2403/A2 U$$882/A1 U$$2403/B2 VGND VGND VPWR VPWR U$$2388/A
+ sky130_fd_sc_hd__a22o_1
XU$$2398 U$$2398/A U$$2442/B VGND VGND VPWR VPWR U$$2398/X sky130_fd_sc_hd__xor2_1
XFILLER_34_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1653 U$$1653/A U$$1679/B VGND VGND VPWR VPWR U$$1653/X sky130_fd_sc_hd__xor2_1
XU$$1664 U$$1799/B1 U$$1696/A2 U$$1666/A1 U$$1696/B2 VGND VGND VPWR VPWR U$$1665/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1675 U$$1675/A U$$1751/B VGND VGND VPWR VPWR U$$1675/X sky130_fd_sc_hd__xor2_1
XFILLER_194_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1686 U$$727/A1 U$$1688/A2 U$$727/B1 U$$1688/B2 VGND VGND VPWR VPWR U$$1687/A sky130_fd_sc_hd__a22o_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1697 U$$1697/A U$$1751/B VGND VGND VPWR VPWR U$$1697/X sky130_fd_sc_hd__xor2_1
XFILLER_203_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4457_1805 VGND VGND VPWR VPWR U$$4457_1805/HI U$$4457/B sky130_fd_sc_hd__conb_1
XFILLER_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_95_1 dadda_fa_5_95_1/A dadda_fa_5_95_1/B dadda_fa_5_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_96_0/B dadda_fa_7_95_0/A sky130_fd_sc_hd__fa_1
XFILLER_116_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_88_0 dadda_fa_5_88_0/A dadda_fa_5_88_0/B dadda_fa_5_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_89_0/A dadda_fa_6_88_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_196_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_751 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$305 final_adder.U$$304/B final_adder.U$$179/X final_adder.U$$177/X
+ VGND VGND VPWR VPWR final_adder.U$$305/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$316 final_adder.U$$318/B final_adder.U$$316/B VGND VGND VPWR VPWR
+ final_adder.U$$442/B sky130_fd_sc_hd__and2_1
XFILLER_84_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater520 U$$340/A2 VGND VGND VPWR VPWR U$$316/A2 sky130_fd_sc_hd__clkbuf_4
Xfinal_adder.U$$327 final_adder.U$$326/B final_adder.U$$201/X final_adder.U$$199/X
+ VGND VGND VPWR VPWR final_adder.U$$327/X sky130_fd_sc_hd__a21o_1
Xrepeater531 U$$2858/A2 VGND VGND VPWR VPWR U$$2868/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$338 final_adder.U$$340/B final_adder.U$$338/B VGND VGND VPWR VPWR
+ final_adder.U$$464/B sky130_fd_sc_hd__and2_1
XTAP_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater542 U$$2711/A2 VGND VGND VPWR VPWR U$$2737/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$349 final_adder.U$$348/B final_adder.U$$223/X final_adder.U$$221/X
+ VGND VGND VPWR VPWR final_adder.U$$349/X sky130_fd_sc_hd__a21o_1
Xrepeater553 U$$2333/X VGND VGND VPWR VPWR U$$2403/A2 sky130_fd_sc_hd__clkbuf_8
Xrepeater564 U$$2316/A2 VGND VGND VPWR VPWR U$$2326/A2 sky130_fd_sc_hd__buf_4
XFILLER_38_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater575 U$$2059/X VGND VGND VPWR VPWR U$$2177/A2 sky130_fd_sc_hd__buf_6
XFILLER_26_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater586 U$$1831/A2 VGND VGND VPWR VPWR U$$1839/A2 sky130_fd_sc_hd__buf_6
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater597 U$$1770/A2 VGND VGND VPWR VPWR U$$1764/A2 sky130_fd_sc_hd__buf_6
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4290 U$$4290/A U$$4294/B VGND VGND VPWR VPWR U$$4290/X sky130_fd_sc_hd__xor2_1
XFILLER_81_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_90_0 dadda_fa_4_90_0/A dadda_fa_4_90_0/B dadda_fa_4_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/A dadda_fa_5_90_1/A sky130_fd_sc_hd__fa_1
XFILLER_88_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_104_2 input134/X dadda_fa_3_104_2/B dadda_fa_3_104_2/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_105_1/A dadda_fa_4_104_2/B sky130_fd_sc_hd__fa_1
XFILLER_135_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_118_0 dadda_fa_6_118_0/A dadda_fa_6_118_0/B dadda_fa_6_118_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_119_0/B dadda_fa_7_118_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$861 final_adder.U$$764/X final_adder.U$$829/X final_adder.U$$765/X
+ VGND VGND VPWR VPWR final_adder.U$$861/X sky130_fd_sc_hd__a21o_2
XU$$700 U$$700/A U$$712/B VGND VGND VPWR VPWR U$$700/X sky130_fd_sc_hd__xor2_1
XFILLER_57_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$711 U$$846/B1 U$$711/A2 U$$711/B1 U$$711/B2 VGND VGND VPWR VPWR U$$712/A sky130_fd_sc_hd__a22o_1
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$883 final_adder.U$$786/X final_adder.U$$619/X final_adder.U$$787/X
+ VGND VGND VPWR VPWR final_adder.U$$883/X sky130_fd_sc_hd__a21o_2
XTAP_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_38_3 dadda_fa_3_38_3/A dadda_fa_3_38_3/B dadda_fa_3_38_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_1/B dadda_fa_4_38_2/CIN sky130_fd_sc_hd__fa_1
XU$$722 U$$722/A U$$740/B VGND VGND VPWR VPWR U$$722/X sky130_fd_sc_hd__xor2_1
XFILLER_44_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$733 U$$733/A1 U$$739/A2 U$$48/B1 U$$739/B2 VGND VGND VPWR VPWR U$$734/A sky130_fd_sc_hd__a22o_1
XFILLER_21_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$744 U$$744/A U$$750/B VGND VGND VPWR VPWR U$$744/X sky130_fd_sc_hd__xor2_1
XFILLER_112_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$755 U$$892/A1 U$$759/A2 U$$757/A1 U$$759/B2 VGND VGND VPWR VPWR U$$756/A sky130_fd_sc_hd__a22o_1
XFILLER_43_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$766 U$$766/A U$$770/B VGND VGND VPWR VPWR U$$766/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$777 U$$914/A1 U$$783/A2 U$$914/B1 U$$783/B2 VGND VGND VPWR VPWR U$$778/A sky130_fd_sc_hd__a22o_1
XFILLER_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$788 U$$788/A U$$794/B VGND VGND VPWR VPWR U$$788/X sky130_fd_sc_hd__xor2_1
XFILLER_71_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$799 U$$799/A1 U$$805/A2 U$$938/A1 U$$805/B2 VGND VGND VPWR VPWR U$$800/A sky130_fd_sc_hd__a22o_1
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1600 U$$4496/A1 VGND VGND VPWR VPWR U$$2715/A1 sky130_fd_sc_hd__buf_4
XFILLER_8_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1611 U$$3944/A1 VGND VGND VPWR VPWR U$$654/B1 sky130_fd_sc_hd__buf_4
XANTENNA_5 _327_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1622 U$$1338/B VGND VGND VPWR VPWR U$$1330/B sky130_fd_sc_hd__buf_6
Xrepeater1633 U$$3987/B1 VGND VGND VPWR VPWR U$$2754/B1 sky130_fd_sc_hd__buf_2
Xrepeater1644 input108/X VGND VGND VPWR VPWR U$$4490/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_99_805 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1655 U$$4484/B1 VGND VGND VPWR VPWR U$$650/A1 sky130_fd_sc_hd__buf_4
Xrepeater1666 U$$3114/A1 VGND VGND VPWR VPWR U$$2701/B1 sky130_fd_sc_hd__buf_6
XFILLER_98_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1677 U$$918/A1 VGND VGND VPWR VPWR U$$916/B1 sky130_fd_sc_hd__buf_6
Xrepeater1688 U$$2834/A1 VGND VGND VPWR VPWR U$$94/A1 sky130_fd_sc_hd__clkbuf_8
Xrepeater1699 U$$3517/A1 VGND VGND VPWR VPWR U$$366/A1 sky130_fd_sc_hd__buf_8
XFILLER_140_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_692 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_40_3 U$$2747/X U$$2755/B input191/X VGND VGND VPWR VPWR dadda_fa_3_41_1/B
+ dadda_fa_3_40_3/B sky130_fd_sc_hd__fa_1
XFILLER_26_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_33_2 U$$871/X U$$1004/X U$$1137/X VGND VGND VPWR VPWR dadda_fa_3_34_1/A
+ dadda_fa_3_33_3/A sky130_fd_sc_hd__fa_1
XFILLER_34_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_10_1 dadda_fa_5_10_1/A dadda_fa_5_10_1/B dadda_ha_4_10_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_11_0/B dadda_fa_7_10_0/A sky130_fd_sc_hd__fa_1
XU$$2140 U$$2140/A U$$2150/B VGND VGND VPWR VPWR U$$2140/X sky130_fd_sc_hd__xor2_1
XFILLER_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2151 U$$918/A1 U$$2189/A2 U$$783/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2152/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_26_1 U$$458/X U$$591/X U$$724/X VGND VGND VPWR VPWR dadda_fa_3_27_2/CIN
+ dadda_fa_3_26_3/CIN sky130_fd_sc_hd__fa_1
XU$$2162 U$$2162/A U$$2184/B VGND VGND VPWR VPWR U$$2162/X sky130_fd_sc_hd__xor2_1
XU$$2173 U$$2445/B1 U$$2177/A2 U$$2312/A1 U$$2177/B2 VGND VGND VPWR VPWR U$$2174/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2184 U$$2184/A U$$2184/B VGND VGND VPWR VPWR U$$2184/X sky130_fd_sc_hd__xor2_1
XU$$1450 U$$4188/B1 U$$1502/A2 U$$4055/A1 U$$1502/B2 VGND VGND VPWR VPWR U$$1451/A
+ sky130_fd_sc_hd__a22o_1
XU$$2195 U$$2311/B U$$2195/B VGND VGND VPWR VPWR U$$2195/X sky130_fd_sc_hd__and2_1
XFILLER_62_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1461 U$$1461/A U$$1506/A VGND VGND VPWR VPWR U$$1461/X sky130_fd_sc_hd__xor2_1
XFILLER_179_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1472 U$$2292/B1 U$$1374/X U$$2842/B1 U$$1375/X VGND VGND VPWR VPWR U$$1473/A sky130_fd_sc_hd__a22o_1
XFILLER_50_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_991 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1483 U$$1483/A U$$1501/B VGND VGND VPWR VPWR U$$1483/X sky130_fd_sc_hd__xor2_1
XU$$1494 U$$946/A1 U$$1502/A2 U$$811/A1 U$$1502/B2 VGND VGND VPWR VPWR U$$1495/A sky130_fd_sc_hd__a22o_1
XFILLER_124_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_85_5 U$$3502/X U$$3635/X U$$3768/X VGND VGND VPWR VPWR dadda_fa_2_86_4/A
+ dadda_fa_3_85_0/A sky130_fd_sc_hd__fa_2
XFILLER_132_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_78_4 U$$2823/X U$$2956/X U$$3089/X VGND VGND VPWR VPWR dadda_fa_2_79_1/CIN
+ dadda_fa_2_78_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_44_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4511_1832 VGND VGND VPWR VPWR U$$4511_1832/HI U$$4511/B sky130_fd_sc_hd__conb_1
XFILLER_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$102 _398_/Q _270_/Q VGND VGND VPWR VPWR final_adder.U$$923/B1 final_adder.U$$152/A
+ sky130_fd_sc_hd__ha_1
XTAP_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$113 _409_/Q _281_/Q VGND VGND VPWR VPWR final_adder.U$$143/B1 final_adder.U$$142/B
+ sky130_fd_sc_hd__ha_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$124 _420_/Q _292_/Q VGND VGND VPWR VPWR final_adder.U$$901/B1 final_adder.U$$130/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_4_48_2 dadda_fa_4_48_2/A dadda_fa_4_48_2/B dadda_fa_4_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/CIN dadda_fa_5_48_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$135 final_adder.U$$134/B final_adder.U$$905/B1 final_adder.U$$135/B1
+ VGND VGND VPWR VPWR final_adder.U$$135/X sky130_fd_sc_hd__a21o_1
XTAP_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$146 final_adder.U$$146/A final_adder.U$$146/B VGND VGND VPWR VPWR
+ final_adder.U$$274/B sky130_fd_sc_hd__and2_1
XTAP_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$157 final_adder.U$$156/B final_adder.U$$927/B1 final_adder.U$$157/B1
+ VGND VGND VPWR VPWR final_adder.U$$157/X sky130_fd_sc_hd__a21o_1
XTAP_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$168 final_adder.U$$168/A final_adder.U$$168/B VGND VGND VPWR VPWR
+ final_adder.U$$296/B sky130_fd_sc_hd__and2_1
XTAP_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$179 final_adder.U$$178/B final_adder.U$$949/B1 final_adder.U$$179/B1
+ VGND VGND VPWR VPWR final_adder.U$$179/X sky130_fd_sc_hd__a21o_1
Xrepeater394 U$$892/A2 VGND VGND VPWR VPWR U$$882/A2 sky130_fd_sc_hd__buf_4
XFILLER_66_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_18_0 dadda_fa_7_18_0/A dadda_fa_7_18_0/B dadda_fa_7_18_0/CIN VGND VGND
+ VPWR VPWR _315_/D _186_/D sky130_fd_sc_hd__fa_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1026 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput120 b[5] VGND VGND VPWR VPWR input120/X sky130_fd_sc_hd__buf_6
XFILLER_209_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput131 c[101] VGND VGND VPWR VPWR input131/X sky130_fd_sc_hd__buf_4
Xdadda_fa_3_50_2 dadda_fa_3_50_2/A dadda_fa_3_50_2/B dadda_fa_3_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_1/A dadda_fa_4_50_2/B sky130_fd_sc_hd__fa_1
Xinput142 c[111] VGND VGND VPWR VPWR input142/X sky130_fd_sc_hd__clkbuf_4
XFILLER_114_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_66_2 U$$937/X U$$1070/X U$$1203/X VGND VGND VPWR VPWR dadda_fa_1_67_6/A
+ dadda_fa_1_66_8/A sky130_fd_sc_hd__fa_1
Xinput153 c[121] VGND VGND VPWR VPWR input153/X sky130_fd_sc_hd__buf_2
XTAP_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput164 c[16] VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__clkbuf_4
XFILLER_114_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 c[26] VGND VGND VPWR VPWR input175/X sky130_fd_sc_hd__clkbuf_2
XTAP_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_43_1 dadda_fa_3_43_1/A dadda_fa_3_43_1/B dadda_fa_3_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_0/CIN dadda_fa_4_43_2/A sky130_fd_sc_hd__fa_1
Xinput186 c[36] VGND VGND VPWR VPWR input186/X sky130_fd_sc_hd__buf_2
XFILLER_91_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_59_1 U$$524/X U$$657/X U$$790/X VGND VGND VPWR VPWR dadda_fa_1_60_6/CIN
+ dadda_fa_1_59_8/B sky130_fd_sc_hd__fa_1
Xinput197 c[46] VGND VGND VPWR VPWR input197/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_20_0 dadda_fa_6_20_0/A dadda_fa_6_20_0/B dadda_fa_6_20_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_21_0/B dadda_fa_7_20_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$680 final_adder.U$$696/B final_adder.U$$680/B VGND VGND VPWR VPWR
+ final_adder.U$$792/B sky130_fd_sc_hd__and2_1
XTAP_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_36_0 dadda_fa_3_36_0/A dadda_fa_3_36_0/B dadda_fa_3_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_0/B dadda_fa_4_36_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$691 final_adder.U$$690/B final_adder.U$$587/X final_adder.U$$571/X
+ VGND VGND VPWR VPWR final_adder.U$$691/X sky130_fd_sc_hd__a21o_1
XTAP_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$530 U$$530/A U$$536/B VGND VGND VPWR VPWR U$$530/X sky130_fd_sc_hd__xor2_1
XTAP_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$541 U$$676/B1 U$$415/X U$$678/B1 U$$416/X VGND VGND VPWR VPWR U$$542/A sky130_fd_sc_hd__a22o_1
XTAP_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$552 U$$550/Y U$$549/A U$$548/A U$$551/X U$$548/Y VGND VGND VPWR VPWR U$$552/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_204_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$563 U$$563/A U$$651/B VGND VGND VPWR VPWR U$$563/X sky130_fd_sc_hd__xor2_1
XTAP_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$574 U$$846/B1 U$$606/A2 U$$850/A1 U$$606/B2 VGND VGND VPWR VPWR U$$575/A sky130_fd_sc_hd__a22o_1
XFILLER_16_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$585 U$$585/A U$$607/B VGND VGND VPWR VPWR U$$585/X sky130_fd_sc_hd__xor2_1
XFILLER_205_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$596 U$$733/A1 U$$616/A2 U$$48/B1 U$$616/B2 VGND VGND VPWR VPWR U$$597/A sky130_fd_sc_hd__a22o_1
XFILLER_204_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_95_4 U$$4187/X U$$4320/X U$$4453/X VGND VGND VPWR VPWR dadda_fa_3_96_1/CIN
+ dadda_fa_3_95_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1430 U$$1779/B VGND VGND VPWR VPWR U$$1739/B sky130_fd_sc_hd__buf_12
Xrepeater1441 U$$1558/B VGND VGND VPWR VPWR U$$1546/B sky130_fd_sc_hd__buf_6
XFILLER_172_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1452 U$$1499/B VGND VGND VPWR VPWR U$$1449/B sky130_fd_sc_hd__buf_6
XFILLER_193_1041 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1463 input128/X VGND VGND VPWR VPWR U$$4408/B1 sky130_fd_sc_hd__buf_4
XFILLER_125_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_88_3 dadda_fa_2_88_3/A dadda_fa_2_88_3/B dadda_fa_2_88_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_1/B dadda_fa_3_88_3/B sky130_fd_sc_hd__fa_1
Xrepeater1474 U$$3447/A1 VGND VGND VPWR VPWR U$$1666/A1 sky130_fd_sc_hd__buf_6
XFILLER_67_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1485 U$$4404/A1 VGND VGND VPWR VPWR U$$3719/A1 sky130_fd_sc_hd__buf_6
Xrepeater1496 input124/X VGND VGND VPWR VPWR U$$3557/B1 sky130_fd_sc_hd__buf_4
XFILLER_114_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_58_1 dadda_fa_5_58_1/A dadda_fa_5_58_1/B dadda_fa_5_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_59_0/B dadda_fa_7_58_0/A sky130_fd_sc_hd__fa_1
XFILLER_80_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_104_1 U$$3141/X U$$3274/X U$$3407/X VGND VGND VPWR VPWR dadda_fa_3_105_3/A
+ dadda_fa_3_104_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1280 U$$1280/A U$$1286/B VGND VGND VPWR VPWR U$$1280/X sky130_fd_sc_hd__xor2_1
XU$$1291 U$$58/A1 U$$1337/A2 U$$60/A1 U$$1291/B2 VGND VGND VPWR VPWR U$$1292/A sky130_fd_sc_hd__a22o_1
XFILLER_195_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_125_0 U$$4246/Y U$$4380/X U$$4513/X VGND VGND VPWR VPWR dadda_fa_6_126_0/CIN
+ dadda_fa_7_125_0/A sky130_fd_sc_hd__fa_1
XFILLER_149_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_23 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_2 U$$2168/X U$$2301/X U$$2434/X VGND VGND VPWR VPWR dadda_fa_2_84_2/B
+ dadda_fa_2_83_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_85_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_60_1 dadda_fa_4_60_1/A dadda_fa_4_60_1/B dadda_fa_4_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/B dadda_fa_5_60_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_76_1 U$$1888/X U$$2021/X U$$2154/X VGND VGND VPWR VPWR dadda_fa_2_77_0/CIN
+ dadda_fa_2_76_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_53_0 dadda_fa_4_53_0/A dadda_fa_4_53_0/B dadda_fa_4_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/A dadda_fa_5_53_1/A sky130_fd_sc_hd__fa_1
XFILLER_131_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_69_0 U$$2406/X U$$2539/X U$$2672/X VGND VGND VPWR VPWR dadda_fa_2_70_0/B
+ dadda_fa_2_69_3/B sky130_fd_sc_hd__fa_1
XFILLER_86_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2909 U$$32/A1 U$$2995/A2 U$$32/B1 U$$2995/B2 VGND VGND VPWR VPWR U$$2910/A sky130_fd_sc_hd__a22o_1
XFILLER_22_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _199_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_225 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 _292_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 U$$4404/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_269 U$$2302/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_590 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_362_ _362_/CLK _362_/D VGND VGND VPWR VPWR _362_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_293_ _422_/CLK _293_/D VGND VGND VPWR VPWR _293_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_195_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_982 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_98_2 dadda_fa_3_98_2/A dadda_fa_3_98_2/B dadda_fa_3_98_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_1/A dadda_fa_4_98_2/B sky130_fd_sc_hd__fa_1
XFILLER_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_86_0_1855 VGND VGND VPWR VPWR dadda_fa_1_86_0/A dadda_fa_1_86_0_1855/LO
+ sky130_fd_sc_hd__conb_1
Xdadda_fa_6_68_0 dadda_fa_6_68_0/A dadda_fa_6_68_0/B dadda_fa_6_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_69_0/B dadda_fa_7_68_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_71_0 U$$547/Y U$$681/X U$$814/X VGND VGND VPWR VPWR dadda_fa_1_72_6/CIN
+ dadda_fa_1_71_8/A sky130_fd_sc_hd__fa_1
XFILLER_111_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_5_7_1 U$$420/X input234/X VGND VGND VPWR VPWR dadda_fa_6_8_0/B dadda_fa_7_7_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$360 U$$86/A1 U$$396/A2 U$$88/A1 U$$396/B2 VGND VGND VPWR VPWR U$$361/A sky130_fd_sc_hd__a22o_1
XFILLER_33_922 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$371 U$$371/A U$$377/B VGND VGND VPWR VPWR U$$371/X sky130_fd_sc_hd__xor2_1
XFILLER_189_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$382 U$$654/B1 U$$394/A2 U$$521/A1 U$$394/B2 VGND VGND VPWR VPWR U$$383/A sky130_fd_sc_hd__a22o_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$393 U$$393/A U$$395/B VGND VGND VPWR VPWR U$$393/X sky130_fd_sc_hd__xor2_1
XFILLER_34_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_93_1 U$$3252/X U$$3385/X U$$3518/X VGND VGND VPWR VPWR dadda_fa_3_94_0/CIN
+ dadda_fa_3_93_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_70_0 dadda_fa_5_70_0/A dadda_fa_5_70_0/B dadda_fa_5_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_71_0/A dadda_fa_6_70_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_86_0 U$$3770/X U$$3903/X U$$4036/X VGND VGND VPWR VPWR dadda_fa_3_87_0/B
+ dadda_fa_3_86_2/B sky130_fd_sc_hd__fa_1
Xrepeater1260 U$$3971/B VGND VGND VPWR VPWR U$$3967/B sky130_fd_sc_hd__buf_6
Xrepeater1271 U$$3836/A VGND VGND VPWR VPWR U$$3778/B sky130_fd_sc_hd__buf_8
Xrepeater1282 U$$959/A VGND VGND VPWR VPWR U$$945/B sky130_fd_sc_hd__buf_6
XFILLER_99_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1293 input49/X VGND VGND VPWR VPWR U$$3643/B sky130_fd_sc_hd__buf_6
Xdadda_ha_1_49_7 U$$2898/X U$$3031/X VGND VGND VPWR VPWR dadda_fa_2_50_3/A dadda_fa_3_49_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_141_584 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_62_7 dadda_fa_1_62_7/A dadda_fa_1_62_7/B dadda_fa_1_62_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_2/CIN dadda_fa_2_62_5/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_1_55_6 U$$3176/X U$$3309/X U$$3442/X VGND VGND VPWR VPWR dadda_fa_2_56_2/B
+ dadda_fa_2_55_5/B sky130_fd_sc_hd__fa_1
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_48_5 U$$2098/X U$$2231/X U$$2364/X VGND VGND VPWR VPWR dadda_fa_2_49_2/CIN
+ dadda_fa_2_48_5/B sky130_fd_sc_hd__fa_1
XFILLER_209_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_7_0 dadda_fa_7_7_0/A dadda_fa_7_7_0/B dadda_fa_7_7_0/CIN VGND VGND VPWR
+ VPWR _304_/D _175_/D sky130_fd_sc_hd__fa_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_85_0 dadda_fa_7_85_0/A dadda_fa_7_85_0/B dadda_fa_7_85_0/CIN VGND VGND
+ VPWR VPWR _382_/D _253_/D sky130_fd_sc_hd__fa_1
XFILLER_128_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_74_0_1850 VGND VGND VPWR VPWR dadda_fa_0_74_0/A dadda_fa_0_74_0_1850/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4108 U$$4108/A input55/X VGND VGND VPWR VPWR U$$4108/X sky130_fd_sc_hd__xor2_1
XU$$4119 U$$4119/A U$$4145/B VGND VGND VPWR VPWR U$$4119/X sky130_fd_sc_hd__xor2_1
XFILLER_58_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3407 U$$3407/A U$$3424/A VGND VGND VPWR VPWR U$$3407/X sky130_fd_sc_hd__xor2_1
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3418 input122/X U$$3422/A2 U$$3555/B1 U$$3422/B2 VGND VGND VPWR VPWR U$$3419/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_100_0 dadda_fa_6_100_0/A dadda_fa_6_100_0/B dadda_fa_6_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_101_0/B dadda_fa_7_100_0/CIN sky130_fd_sc_hd__fa_1
XU$$3429 U$$3427/Y input46/X U$$3377/B U$$3428/X U$$3425/Y VGND VGND VPWR VPWR U$$3429/X
+ sky130_fd_sc_hd__a32o_4
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2706 U$$2706/A U$$2710/B VGND VGND VPWR VPWR U$$2706/X sky130_fd_sc_hd__xor2_1
XFILLER_46_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2717 U$$2717/A1 U$$2737/A2 U$$4361/B1 U$$2737/B2 VGND VGND VPWR VPWR U$$2718/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2728 U$$2728/A U$$2736/B VGND VGND VPWR VPWR U$$2728/X sky130_fd_sc_hd__xor2_1
XFILLER_34_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2739 U$$2739/A VGND VGND VPWR VPWR U$$2739/Y sky130_fd_sc_hd__inv_1
XFILLER_61_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1032 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ _414_/CLK _414_/D VGND VGND VPWR VPWR _414_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ _345_/CLK _345_/D VGND VGND VPWR VPWR _345_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_144_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_276_ _407_/CLK _276_/D VGND VGND VPWR VPWR _276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_668 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_65_5 dadda_fa_2_65_5/A dadda_fa_2_65_5/B dadda_fa_2_65_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_2/A dadda_fa_4_65_0/A sky130_fd_sc_hd__fa_2
XFILLER_97_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater905 U$$2415/B1 VGND VGND VPWR VPWR U$$88/A1 sky130_fd_sc_hd__buf_4
XFILLER_68_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater916 input98/X VGND VGND VPWR VPWR U$$4398/A1 sky130_fd_sc_hd__clkbuf_8
Xrepeater927 U$$4055/B1 VGND VGND VPWR VPWR U$$84/A1 sky130_fd_sc_hd__buf_6
Xrepeater938 U$$2409/B1 VGND VGND VPWR VPWR U$$630/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_58_4 dadda_fa_2_58_4/A dadda_fa_2_58_4/B dadda_fa_2_58_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/CIN dadda_fa_3_58_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater949 input94/X VGND VGND VPWR VPWR U$$3642/A1 sky130_fd_sc_hd__buf_6
XFILLER_37_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3930 U$$4476/B1 U$$3946/A2 U$$4343/A1 U$$3946/B2 VGND VGND VPWR VPWR U$$3931/A
+ sky130_fd_sc_hd__a22o_1
XU$$3941 U$$3941/A U$$3967/B VGND VGND VPWR VPWR U$$3941/X sky130_fd_sc_hd__xor2_1
XFILLER_92_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3952 input114/X U$$3968/A2 input115/X U$$3968/B2 VGND VGND VPWR VPWR U$$3953/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3963 U$$3963/A U$$3967/B VGND VGND VPWR VPWR U$$3963/X sky130_fd_sc_hd__xor2_1
XFILLER_80_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3974 input54/X VGND VGND VPWR VPWR U$$3976/B sky130_fd_sc_hd__inv_1
XU$$3985 U$$4396/A1 U$$4011/A2 U$$4398/A1 U$$4011/B2 VGND VGND VPWR VPWR U$$3986/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3996 U$$3996/A U$$4036/B VGND VGND VPWR VPWR U$$3996/X sky130_fd_sc_hd__xor2_1
XFILLER_17_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$190 U$$190/A U$$218/B VGND VGND VPWR VPWR U$$190/X sky130_fd_sc_hd__xor2_1
XFILLER_178_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_941 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput265 output265/A VGND VGND VPWR VPWR o[107] sky130_fd_sc_hd__buf_2
Xoutput276 output276/A VGND VGND VPWR VPWR o[117] sky130_fd_sc_hd__buf_2
XFILLER_47_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1090 U$$3473/A1 VGND VGND VPWR VPWR U$$594/B1 sky130_fd_sc_hd__buf_8
XFILLER_88_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput287 output287/A VGND VGND VPWR VPWR o[127] sky130_fd_sc_hd__buf_2
XFILLER_82_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput298 output298/A VGND VGND VPWR VPWR o[21] sky130_fd_sc_hd__buf_2
XFILLER_181_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_60_4 U$$3585/X U$$3718/X U$$3851/X VGND VGND VPWR VPWR dadda_fa_2_61_1/CIN
+ dadda_fa_2_60_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_53_3 U$$1576/X U$$1709/X U$$1842/X VGND VGND VPWR VPWR dadda_fa_2_54_1/B
+ dadda_fa_2_53_4/B sky130_fd_sc_hd__fa_1
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_30_2 dadda_fa_4_30_2/A dadda_fa_4_30_2/B dadda_fa_4_30_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/CIN dadda_fa_5_30_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_46_2 U$$897/X U$$1030/X U$$1163/X VGND VGND VPWR VPWR dadda_fa_2_47_2/B
+ dadda_fa_2_46_4/CIN sky130_fd_sc_hd__fa_2
XFILLER_16_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_23_1 dadda_fa_4_23_1/A dadda_fa_4_23_1/B dadda_fa_4_23_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/B dadda_fa_5_23_1/B sky130_fd_sc_hd__fa_1
XFILLER_167_1046 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_39_1 U$$484/X U$$617/X U$$750/X VGND VGND VPWR VPWR dadda_fa_2_40_4/B
+ dadda_fa_2_39_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_16_0 U$$704/X U$$837/X U$$970/X VGND VGND VPWR VPWR dadda_fa_5_17_0/A
+ dadda_fa_5_16_1/A sky130_fd_sc_hd__fa_1
XFILLER_130_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1106 final_adder.U$$172/A final_adder.U$$881/X VGND VGND VPWR VPWR
+ output365/A sky130_fd_sc_hd__xor2_1
XFILLER_184_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1117 final_adder.U$$162/B final_adder.U$$933/X VGND VGND VPWR VPWR
+ output377/A sky130_fd_sc_hd__xor2_1
XFILLER_149_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1128 final_adder.U$$150/A final_adder.U$$859/X VGND VGND VPWR VPWR
+ output262/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1139 final_adder.U$$140/B final_adder.U$$911/X VGND VGND VPWR VPWR
+ output274/A sky130_fd_sc_hd__xor2_1
XFILLER_183_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1036 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_68_3 dadda_fa_3_68_3/A dadda_fa_3_68_3/B dadda_fa_3_68_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_1/B dadda_fa_4_68_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3204 U$$3204/A U$$3242/B VGND VGND VPWR VPWR U$$3204/X sky130_fd_sc_hd__xor2_1
XFILLER_59_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3215 U$$3215/A1 U$$3229/A2 U$$4450/A1 U$$3227/B2 VGND VGND VPWR VPWR U$$3216/A
+ sky130_fd_sc_hd__a22o_1
XU$$3226 U$$3226/A U$$3288/A VGND VGND VPWR VPWR U$$3226/X sky130_fd_sc_hd__xor2_1
XFILLER_207_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$19 _315_/Q _187_/Q VGND VGND VPWR VPWR final_adder.U$$237/B1 final_adder.U$$236/B
+ sky130_fd_sc_hd__ha_1
XU$$3237 U$$3511/A1 U$$3241/A2 U$$3376/A1 U$$3241/B2 VGND VGND VPWR VPWR U$$3238/A
+ sky130_fd_sc_hd__a22o_1
XU$$3248 U$$3248/A U$$3256/B VGND VGND VPWR VPWR U$$3248/X sky130_fd_sc_hd__xor2_1
XU$$2503 U$$2503/A U$$2597/B VGND VGND VPWR VPWR U$$2503/X sky130_fd_sc_hd__xor2_1
XU$$3259 U$$654/B1 U$$3263/A2 U$$521/A1 U$$3263/B2 VGND VGND VPWR VPWR U$$3260/A sky130_fd_sc_hd__a22o_1
XU$$2514 U$$3882/B1 U$$2600/A2 U$$3749/A1 U$$2600/B2 VGND VGND VPWR VPWR U$$2515/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2525 U$$2525/A U$$2525/B VGND VGND VPWR VPWR U$$2525/X sky130_fd_sc_hd__xor2_1
XFILLER_62_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2536 U$$2808/B1 U$$2558/A2 U$$894/A1 U$$2558/B2 VGND VGND VPWR VPWR U$$2537/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2547 U$$2547/A U$$2569/B VGND VGND VPWR VPWR U$$2547/X sky130_fd_sc_hd__xor2_1
XU$$1802 U$$1802/A U$$1840/B VGND VGND VPWR VPWR U$$1802/X sky130_fd_sc_hd__xor2_1
XU$$1813 U$$991/A1 U$$1819/A2 U$$993/A1 U$$1819/B2 VGND VGND VPWR VPWR U$$1814/A sky130_fd_sc_hd__a22o_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2558 U$$366/A1 U$$2558/A2 U$$2834/A1 U$$2558/B2 VGND VGND VPWR VPWR U$$2559/A
+ sky130_fd_sc_hd__a22o_1
XU$$1824 U$$1824/A U$$1870/B VGND VGND VPWR VPWR U$$1824/X sky130_fd_sc_hd__xor2_1
XU$$2569 U$$2569/A U$$2569/B VGND VGND VPWR VPWR U$$2569/X sky130_fd_sc_hd__xor2_1
XFILLER_62_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1835 U$$52/B1 U$$1839/A2 U$$3481/A1 U$$1839/B2 VGND VGND VPWR VPWR U$$1836/A sky130_fd_sc_hd__a22o_1
XU$$1846 U$$1846/A U$$1880/B VGND VGND VPWR VPWR U$$1846/X sky130_fd_sc_hd__xor2_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1857 U$$759/B1 U$$1869/A2 U$$3366/A1 U$$1869/B2 VGND VGND VPWR VPWR U$$1858/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1868 U$$1868/A U$$1870/B VGND VGND VPWR VPWR U$$1868/X sky130_fd_sc_hd__xor2_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1879 U$$2016/A1 U$$1879/A2 U$$98/B1 U$$1879/B2 VGND VGND VPWR VPWR U$$1880/A sky130_fd_sc_hd__a22o_1
XFILLER_187_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_396 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_328_ _329_/CLK _328_/D VGND VGND VPWR VPWR _328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_259_ _421_/CLK _259_/D VGND VGND VPWR VPWR _259_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_1046 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$554_1838 VGND VGND VPWR VPWR U$$554_1838/HI U$$554/A1 sky130_fd_sc_hd__conb_1
XFILLER_171_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_70_3 dadda_fa_2_70_3/A dadda_fa_2_70_3/B dadda_fa_2_70_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/B dadda_fa_3_70_3/B sky130_fd_sc_hd__fa_1
XFILLER_96_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_63_2 dadda_fa_2_63_2/A dadda_fa_2_63_2/B dadda_fa_2_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/A dadda_fa_3_63_3/A sky130_fd_sc_hd__fa_1
XFILLER_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater702 U$$3874/B2 VGND VGND VPWR VPWR U$$3878/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$509 final_adder.U$$508/B final_adder.U$$393/X final_adder.U$$385/X
+ VGND VGND VPWR VPWR final_adder.U$$509/X sky130_fd_sc_hd__a21o_1
Xrepeater713 U$$3833/B2 VGND VGND VPWR VPWR U$$3819/B2 sky130_fd_sc_hd__buf_6
XFILLER_84_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_40_1 dadda_fa_5_40_1/A dadda_fa_5_40_1/B dadda_fa_5_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_41_0/B dadda_fa_7_40_0/A sky130_fd_sc_hd__fa_2
XFILLER_84_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater724 U$$3567/X VGND VGND VPWR VPWR U$$3644/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_56_1 dadda_fa_2_56_1/A dadda_fa_2_56_1/B dadda_fa_2_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_0/CIN dadda_fa_3_56_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater735 U$$3346/B2 VGND VGND VPWR VPWR U$$3320/B2 sky130_fd_sc_hd__buf_6
Xrepeater746 U$$3255/B2 VGND VGND VPWR VPWR U$$3263/B2 sky130_fd_sc_hd__buf_4
Xrepeater757 U$$3019/X VGND VGND VPWR VPWR U$$3118/B2 sky130_fd_sc_hd__buf_8
Xdadda_fa_5_33_0 dadda_fa_5_33_0/A dadda_fa_5_33_0/B dadda_fa_5_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_34_0/A dadda_fa_6_33_0/CIN sky130_fd_sc_hd__fa_1
XU$$4450 U$$4450/A1 U$$4388/X U$$4452/A1 U$$4476/B2 VGND VGND VPWR VPWR U$$4451/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater768 U$$340/B2 VGND VGND VPWR VPWR U$$302/B2 sky130_fd_sc_hd__buf_4
XFILLER_42_1175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4461 U$$4461/A U$$4461/B VGND VGND VPWR VPWR U$$4461/X sky130_fd_sc_hd__xor2_1
Xrepeater779 U$$2874/B2 VGND VGND VPWR VPWR U$$2858/B2 sky130_fd_sc_hd__buf_4
XFILLER_38_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_49_0 U$$3164/X U$$3297/X input200/X VGND VGND VPWR VPWR dadda_fa_3_50_0/B
+ dadda_fa_3_49_2/B sky130_fd_sc_hd__fa_1
XU$$4472 input99/X U$$4388/X input100/X U$$4486/B2 VGND VGND VPWR VPWR U$$4473/A sky130_fd_sc_hd__a22o_1
XU$$4483 U$$4483/A U$$4483/B VGND VGND VPWR VPWR U$$4483/X sky130_fd_sc_hd__xor2_1
XFILLER_25_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4494 U$$4494/A1 U$$4388/X U$$4496/A1 U$$4494/B2 VGND VGND VPWR VPWR U$$4495/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3760 U$$3760/A U$$3778/B VGND VGND VPWR VPWR U$$3760/X sky130_fd_sc_hd__xor2_1
XU$$3771 U$$4043/B1 U$$3773/A2 U$$3908/B1 U$$3773/B2 VGND VGND VPWR VPWR U$$3772/A
+ sky130_fd_sc_hd__a22o_1
XU$$3782 U$$3782/A U$$3834/B VGND VGND VPWR VPWR U$$3782/X sky130_fd_sc_hd__xor2_1
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3793 U$$4476/B1 U$$3793/A2 U$$4343/A1 U$$3793/B2 VGND VGND VPWR VPWR U$$3794/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_579 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_78_2 dadda_fa_4_78_2/A dadda_fa_4_78_2/B dadda_fa_4_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/CIN dadda_fa_5_78_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_48_0 dadda_fa_7_48_0/A dadda_fa_7_48_0/B dadda_fa_7_48_0/CIN VGND VGND
+ VPWR VPWR _345_/D _216_/D sky130_fd_sc_hd__fa_1
XFILLER_134_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_980 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_96_0_1872 VGND VGND VPWR VPWR dadda_ha_1_96_0/A dadda_ha_1_96_0_1872/LO
+ sky130_fd_sc_hd__conb_1
Xdadda_fa_1_51_0 U$$109/X U$$242/X U$$375/X VGND VGND VPWR VPWR dadda_fa_2_52_0/B
+ dadda_fa_2_51_3/B sky130_fd_sc_hd__fa_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$904 U$$82/A1 U$$906/A2 U$$84/A1 U$$906/B2 VGND VGND VPWR VPWR U$$905/A sky130_fd_sc_hd__a22o_1
XU$$915 U$$915/A U$$919/B VGND VGND VPWR VPWR U$$915/X sky130_fd_sc_hd__xor2_1
XFILLER_141_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$926 U$$926/A1 U$$938/A2 U$$928/A1 U$$938/B2 VGND VGND VPWR VPWR U$$927/A sky130_fd_sc_hd__a22o_1
XU$$937 U$$937/A U$$959/A VGND VGND VPWR VPWR U$$937/X sky130_fd_sc_hd__xor2_1
XFILLER_55_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$948 U$$948/A1 U$$826/X U$$950/A1 U$$827/X VGND VGND VPWR VPWR U$$949/A sky130_fd_sc_hd__a22o_1
XFILLER_83_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$959 U$$959/A VGND VGND VPWR VPWR U$$959/Y sky130_fd_sc_hd__inv_1
XFILLER_55_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1109 U$$1109/A U$$1139/B VGND VGND VPWR VPWR U$$1109/X sky130_fd_sc_hd__xor2_1
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_532 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1057 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_80_2 dadda_fa_3_80_2/A dadda_fa_3_80_2/B dadda_fa_3_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_1/A dadda_fa_4_80_2/B sky130_fd_sc_hd__fa_1
XFILLER_125_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_73_1 dadda_fa_3_73_1/A dadda_fa_3_73_1/B dadda_fa_3_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_0/CIN dadda_fa_4_73_2/A sky130_fd_sc_hd__fa_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_50_0 dadda_fa_6_50_0/A dadda_fa_6_50_0/B dadda_fa_6_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_51_0/B dadda_fa_7_50_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_66_0 dadda_fa_3_66_0/A dadda_fa_3_66_0/B dadda_fa_3_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_0/B dadda_fa_4_66_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_310 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3001 U$$3547/B1 U$$3011/A2 U$$3414/A1 U$$3011/B2 VGND VGND VPWR VPWR U$$3002/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_clk _219_/CLK VGND VGND VPWR VPWR _345_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3012 U$$3012/A U$$3013/A VGND VGND VPWR VPWR U$$3012/X sky130_fd_sc_hd__xor2_1
XFILLER_75_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3023 U$$3023/A U$$3075/B VGND VGND VPWR VPWR U$$3023/X sky130_fd_sc_hd__xor2_1
XU$$3034 U$$4404/A1 U$$3082/A2 U$$981/A1 U$$3082/B2 VGND VGND VPWR VPWR U$$3035/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3045 U$$3045/A U$$3125/B VGND VGND VPWR VPWR U$$3045/X sky130_fd_sc_hd__xor2_1
XU$$2300 U$$2848/A1 U$$2316/A2 U$$2711/B1 U$$2316/B2 VGND VGND VPWR VPWR U$$2301/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2311 U$$2311/A U$$2311/B VGND VGND VPWR VPWR U$$2311/X sky130_fd_sc_hd__xor2_1
XFILLER_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3056 U$$3876/B1 U$$3060/A2 U$$3058/A1 U$$3060/B2 VGND VGND VPWR VPWR U$$3057/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_102_1 dadda_fa_4_102_1/A dadda_fa_4_102_1/B dadda_fa_4_102_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/B dadda_fa_5_102_1/B sky130_fd_sc_hd__fa_1
XFILLER_35_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2322 U$$952/A1 U$$2326/A2 U$$2324/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2323/A
+ sky130_fd_sc_hd__a22o_1
XU$$3067 U$$3067/A U$$3109/B VGND VGND VPWR VPWR U$$3067/X sky130_fd_sc_hd__xor2_1
XU$$2333 U$$2331/Y input28/X input27/X U$$2332/X U$$2329/Y VGND VGND VPWR VPWR U$$2333/X
+ sky130_fd_sc_hd__a32o_4
XU$$3078 U$$3352/A1 U$$3082/A2 U$$3078/B1 U$$3082/B2 VGND VGND VPWR VPWR U$$3079/A
+ sky130_fd_sc_hd__a22o_1
XU$$3089 U$$3089/A U$$3117/B VGND VGND VPWR VPWR U$$3089/X sky130_fd_sc_hd__xor2_1
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2344 U$$2344/A U$$2360/B VGND VGND VPWR VPWR U$$2344/X sky130_fd_sc_hd__xor2_1
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2355 U$$2492/A1 U$$2359/A2 U$$3453/A1 U$$2359/B2 VGND VGND VPWR VPWR U$$2356/A
+ sky130_fd_sc_hd__a22o_1
XU$$1610 U$$1610/A U$$1628/B VGND VGND VPWR VPWR U$$1610/X sky130_fd_sc_hd__xor2_1
XU$$1621 U$$660/B1 U$$1621/A2 U$$388/B1 U$$1621/B2 VGND VGND VPWR VPWR U$$1622/A sky130_fd_sc_hd__a22o_1
XU$$2366 U$$2366/A U$$2366/B VGND VGND VPWR VPWR U$$2366/X sky130_fd_sc_hd__xor2_1
XU$$1632 U$$1632/A U$$1638/B VGND VGND VPWR VPWR U$$1632/X sky130_fd_sc_hd__xor2_1
XU$$2377 U$$3882/B1 U$$2463/A2 U$$3749/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2378/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1643 U$$1644/A VGND VGND VPWR VPWR U$$1643/Y sky130_fd_sc_hd__inv_1
XU$$2388 U$$2388/A U$$2426/B VGND VGND VPWR VPWR U$$2388/X sky130_fd_sc_hd__xor2_1
XFILLER_201_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2399 U$$2808/B1 U$$2333/X U$$894/A1 U$$2334/X VGND VGND VPWR VPWR U$$2400/A sky130_fd_sc_hd__a22o_1
XFILLER_37_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1654 U$$2063/B1 U$$1688/A2 U$$2065/B1 U$$1688/B2 VGND VGND VPWR VPWR U$$1655/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1665 U$$1665/A U$$1679/B VGND VGND VPWR VPWR U$$1665/X sky130_fd_sc_hd__xor2_1
XFILLER_203_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1676 U$$991/A1 U$$1696/A2 U$$2363/A1 U$$1696/B2 VGND VGND VPWR VPWR U$$1677/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1687 U$$1687/A U$$1689/B VGND VGND VPWR VPWR U$$1687/X sky130_fd_sc_hd__xor2_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_123_0 dadda_fa_7_123_0/A dadda_fa_7_123_0/B dadda_fa_7_123_0/CIN VGND
+ VGND VPWR VPWR _420_/D _291_/D sky130_fd_sc_hd__fa_2
XFILLER_188_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1698 U$$874/B1 U$$1706/A2 U$$741/A1 U$$1706/B2 VGND VGND VPWR VPWR U$$1699/A sky130_fd_sc_hd__a22o_1
XFILLER_187_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_88_1 dadda_fa_5_88_1/A dadda_fa_5_88_1/B dadda_fa_5_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_89_0/B dadda_fa_7_88_0/A sky130_fd_sc_hd__fa_2
XFILLER_143_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$306 final_adder.U$$308/B final_adder.U$$306/B VGND VGND VPWR VPWR
+ final_adder.U$$432/B sky130_fd_sc_hd__and2_1
Xrepeater510 U$$3018/X VGND VGND VPWR VPWR U$$3118/A2 sky130_fd_sc_hd__buf_8
Xfinal_adder.U$$317 final_adder.U$$316/B final_adder.U$$191/X final_adder.U$$189/X
+ VGND VGND VPWR VPWR final_adder.U$$317/X sky130_fd_sc_hd__a21o_1
Xrepeater521 U$$340/A2 VGND VGND VPWR VPWR U$$302/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$328 final_adder.U$$330/B final_adder.U$$328/B VGND VGND VPWR VPWR
+ final_adder.U$$454/B sky130_fd_sc_hd__and2_1
Xrepeater532 U$$2874/A2 VGND VGND VPWR VPWR U$$2858/A2 sky130_fd_sc_hd__buf_4
XFILLER_211_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$339 final_adder.U$$338/B final_adder.U$$213/X final_adder.U$$211/X
+ VGND VGND VPWR VPWR final_adder.U$$339/X sky130_fd_sc_hd__a21o_1
XFILLER_57_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater543 U$$2607/X VGND VGND VPWR VPWR U$$2711/A2 sky130_fd_sc_hd__buf_6
XFILLER_38_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_49_clk _239_/CLK VGND VGND VPWR VPWR _367_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_73_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater554 U$$2435/A2 VGND VGND VPWR VPWR U$$2417/A2 sky130_fd_sc_hd__buf_6
Xrepeater565 U$$2196/X VGND VGND VPWR VPWR U$$2316/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_66_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater576 U$$1990/A2 VGND VGND VPWR VPWR U$$1970/A2 sky130_fd_sc_hd__buf_6
XFILLER_37_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater587 U$$1879/A2 VGND VGND VPWR VPWR U$$1831/A2 sky130_fd_sc_hd__buf_8
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4280 U$$4280/A U$$4330/B VGND VGND VPWR VPWR U$$4280/X sky130_fd_sc_hd__xor2_1
XFILLER_26_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater598 U$$1770/A2 VGND VGND VPWR VPWR U$$1746/A2 sky130_fd_sc_hd__buf_8
XFILLER_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4291 U$$4428/A1 U$$4297/A2 U$$4430/A1 U$$4297/B2 VGND VGND VPWR VPWR U$$4292/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3590 U$$4275/A1 U$$3606/A2 U$$3727/B1 U$$3606/B2 VGND VGND VPWR VPWR U$$3591/A
+ sky130_fd_sc_hd__a22o_1
XU$$4505_1829 VGND VGND VPWR VPWR U$$4505_1829/HI U$$4505/B sky130_fd_sc_hd__conb_1
XFILLER_25_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4397_1775 VGND VGND VPWR VPWR U$$4397_1775/HI U$$4397/B sky130_fd_sc_hd__conb_1
Xdadda_fa_4_90_1 dadda_fa_4_90_1/A dadda_fa_4_90_1/B dadda_fa_4_90_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/B dadda_fa_5_90_1/B sky130_fd_sc_hd__fa_1
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_398 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_83_0 dadda_fa_4_83_0/A dadda_fa_4_83_0/B dadda_fa_4_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/A dadda_fa_5_83_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_104_3 dadda_fa_3_104_3/A dadda_fa_3_104_3/B dadda_fa_3_104_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_105_1/B dadda_fa_4_104_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$851 final_adder.U$$754/X final_adder.U$$819/X final_adder.U$$755/X
+ VGND VGND VPWR VPWR final_adder.U$$851/X sky130_fd_sc_hd__a21o_2
XTAP_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$701 U$$975/A1 U$$711/A2 U$$703/A1 U$$711/B2 VGND VGND VPWR VPWR U$$702/A sky130_fd_sc_hd__a22o_1
XFILLER_91_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$873 final_adder.U$$776/X final_adder.U$$729/X final_adder.U$$777/X
+ VGND VGND VPWR VPWR ANTENNA_250/DIODE sky130_fd_sc_hd__a21o_1
XTAP_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$712 U$$712/A U$$712/B VGND VGND VPWR VPWR U$$712/X sky130_fd_sc_hd__xor2_1
XU$$723 U$$860/A1 U$$759/A2 U$$860/B1 U$$759/B2 VGND VGND VPWR VPWR U$$724/A sky130_fd_sc_hd__a22o_1
XFILLER_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$895 final_adder.U$$798/X final_adder.U$$381/X final_adder.U$$799/X
+ VGND VGND VPWR VPWR final_adder.U$$895/X sky130_fd_sc_hd__a21o_1
XFILLER_17_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$734 U$$734/A U$$740/B VGND VGND VPWR VPWR U$$734/X sky130_fd_sc_hd__xor2_1
XU$$745 U$$745/A1 U$$749/A2 U$$882/B1 U$$749/B2 VGND VGND VPWR VPWR U$$746/A sky130_fd_sc_hd__a22o_1
XFILLER_21_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$756 U$$756/A U$$796/B VGND VGND VPWR VPWR U$$756/X sky130_fd_sc_hd__xor2_1
XFILLER_205_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$767 U$$82/A1 U$$793/A2 U$$84/A1 U$$793/B2 VGND VGND VPWR VPWR U$$768/A sky130_fd_sc_hd__a22o_1
XFILLER_189_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$778 U$$778/A U$$784/B VGND VGND VPWR VPWR U$$778/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$789 U$$789/A1 U$$689/X U$$928/A1 U$$690/X VGND VGND VPWR VPWR U$$790/A sky130_fd_sc_hd__a22o_1
Xclkbuf_3_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _219_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_204_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_98_0 dadda_fa_6_98_0/A dadda_fa_6_98_0/B dadda_fa_6_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_99_0/B dadda_fa_7_98_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1601 U$$4496/A1 VGND VGND VPWR VPWR U$$521/B1 sky130_fd_sc_hd__buf_6
XANTENNA_6 _327_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1612 U$$2848/A1 VGND VGND VPWR VPWR U$$2709/B1 sky130_fd_sc_hd__buf_4
XFILLER_137_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1623 U$$1370/A VGND VGND VPWR VPWR U$$1338/B sky130_fd_sc_hd__buf_8
Xrepeater1634 U$$3987/B1 VGND VGND VPWR VPWR U$$4400/A1 sky130_fd_sc_hd__buf_6
Xrepeater1645 U$$652/A1 VGND VGND VPWR VPWR U$$926/A1 sky130_fd_sc_hd__buf_6
Xrepeater1656 U$$2292/B1 VGND VGND VPWR VPWR U$$2842/A1 sky130_fd_sc_hd__buf_4
XFILLER_99_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1667 U$$4484/A1 VGND VGND VPWR VPWR U$$3114/A1 sky130_fd_sc_hd__buf_6
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1678 U$$4478/B1 VGND VGND VPWR VPWR U$$918/A1 sky130_fd_sc_hd__clkbuf_8
Xrepeater1689 U$$2834/A1 VGND VGND VPWR VPWR U$$3108/A1 sky130_fd_sc_hd__buf_6
XFILLER_113_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_40_4 dadda_fa_2_40_4/A dadda_fa_2_40_4/B dadda_fa_2_40_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_41_1/CIN dadda_fa_3_40_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_33_3 U$$1270/X U$$1403/X U$$1536/X VGND VGND VPWR VPWR dadda_fa_3_34_1/B
+ dadda_fa_3_33_3/B sky130_fd_sc_hd__fa_1
XU$$2130 U$$2130/A U$$2170/B VGND VGND VPWR VPWR U$$2130/X sky130_fd_sc_hd__xor2_1
XFILLER_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2141 U$$3235/B1 U$$2169/A2 U$$2691/A1 U$$2169/B2 VGND VGND VPWR VPWR U$$2142/A
+ sky130_fd_sc_hd__a22o_1
XU$$2152 U$$2152/A U$$2191/A VGND VGND VPWR VPWR U$$2152/X sky130_fd_sc_hd__xor2_1
XU$$2163 U$$2848/A1 U$$2183/A2 U$$2165/A1 U$$2183/B2 VGND VGND VPWR VPWR U$$2164/A
+ sky130_fd_sc_hd__a22o_1
XU$$2174 U$$2174/A U$$2178/B VGND VGND VPWR VPWR U$$2174/X sky130_fd_sc_hd__xor2_1
XU$$2185 U$$3829/A1 U$$2189/A2 U$$4103/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2186/A
+ sky130_fd_sc_hd__a22o_1
XU$$1440 U$$1714/A1 U$$1448/A2 U$$72/A1 U$$1448/B2 VGND VGND VPWR VPWR U$$1441/A sky130_fd_sc_hd__a22o_1
XFILLER_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1451 U$$1451/A U$$1499/B VGND VGND VPWR VPWR U$$1451/X sky130_fd_sc_hd__xor2_1
XU$$2196 U$$2194/Y input26/X input25/X U$$2195/X U$$2192/Y VGND VGND VPWR VPWR U$$2196/X
+ sky130_fd_sc_hd__a32o_4
XU$$1462 U$$92/A1 U$$1462/A2 U$$94/A1 U$$1462/B2 VGND VGND VPWR VPWR U$$1463/A sky130_fd_sc_hd__a22o_1
XU$$1473 U$$1473/A U$$1507/A VGND VGND VPWR VPWR U$$1473/X sky130_fd_sc_hd__xor2_1
XFILLER_50_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1484 U$$2717/A1 U$$1504/A2 U$$527/A1 U$$1504/B2 VGND VGND VPWR VPWR U$$1485/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1495 U$$1495/A U$$1499/B VGND VGND VPWR VPWR U$$1495/X sky130_fd_sc_hd__xor2_1
XFILLER_30_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_78_5 U$$3222/X U$$3355/X U$$3488/X VGND VGND VPWR VPWR dadda_fa_2_79_2/A
+ dadda_fa_2_78_5/A sky130_fd_sc_hd__fa_1
XFILLER_44_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$103 _399_/Q _271_/Q VGND VGND VPWR VPWR final_adder.U$$153/B1 final_adder.U$$152/B
+ sky130_fd_sc_hd__ha_1
XTAP_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$114 _410_/Q _282_/Q VGND VGND VPWR VPWR final_adder.U$$911/B1 final_adder.U$$140/A
+ sky130_fd_sc_hd__ha_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$125 _421_/Q _293_/Q VGND VGND VPWR VPWR final_adder.U$$131/B1 final_adder.U$$130/B
+ sky130_fd_sc_hd__ha_1
XFILLER_111_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$136 final_adder.U$$136/A final_adder.U$$136/B VGND VGND VPWR VPWR
+ final_adder.U$$264/B sky130_fd_sc_hd__and2_1
XTAP_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$147 final_adder.U$$146/B final_adder.U$$917/B1 final_adder.U$$147/B1
+ VGND VGND VPWR VPWR final_adder.U$$147/X sky130_fd_sc_hd__a21o_1
XTAP_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$158 final_adder.U$$158/A final_adder.U$$158/B VGND VGND VPWR VPWR
+ final_adder.U$$286/B sky130_fd_sc_hd__and2_1
XTAP_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$169 final_adder.U$$168/B final_adder.U$$939/B1 final_adder.U$$169/B1
+ VGND VGND VPWR VPWR final_adder.U$$169/X sky130_fd_sc_hd__a21o_2
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater395 U$$938/A2 VGND VGND VPWR VPWR U$$892/A2 sky130_fd_sc_hd__buf_6
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1038 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_102_0 U$$4068/X U$$4201/X U$$4334/X VGND VGND VPWR VPWR dadda_fa_4_103_0/B
+ dadda_fa_4_102_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_107_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput110 b[50] VGND VGND VPWR VPWR input110/X sky130_fd_sc_hd__buf_6
XFILLER_88_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput121 b[60] VGND VGND VPWR VPWR input121/X sky130_fd_sc_hd__buf_6
XFILLER_62_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput132 c[102] VGND VGND VPWR VPWR input132/X sky130_fd_sc_hd__buf_4
XFILLER_209_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput143 c[112] VGND VGND VPWR VPWR input143/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_50_3 dadda_fa_3_50_3/A dadda_fa_3_50_3/B dadda_fa_3_50_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_1/B dadda_fa_4_50_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_66_3 U$$1336/X U$$1469/X U$$1602/X VGND VGND VPWR VPWR dadda_fa_1_67_6/B
+ dadda_fa_1_66_8/B sky130_fd_sc_hd__fa_1
Xinput154 c[122] VGND VGND VPWR VPWR input154/X sky130_fd_sc_hd__buf_2
XFILLER_49_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput165 c[17] VGND VGND VPWR VPWR input165/X sky130_fd_sc_hd__clkbuf_4
XTAP_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_43_2 dadda_fa_3_43_2/A dadda_fa_3_43_2/B dadda_fa_3_43_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_1/A dadda_fa_4_43_2/B sky130_fd_sc_hd__fa_1
Xinput176 c[27] VGND VGND VPWR VPWR input176/X sky130_fd_sc_hd__clkbuf_2
XTAP_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput187 c[37] VGND VGND VPWR VPWR input187/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput198 c[47] VGND VGND VPWR VPWR input198/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_0_59_2 U$$923/X U$$1056/X U$$1189/X VGND VGND VPWR VPWR dadda_fa_1_60_7/A
+ dadda_fa_1_59_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$670 final_adder.U$$686/B final_adder.U$$670/B VGND VGND VPWR VPWR
+ final_adder.U$$782/B sky130_fd_sc_hd__and2_1
XTAP_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$681 final_adder.U$$680/B final_adder.U$$577/X final_adder.U$$561/X
+ VGND VGND VPWR VPWR final_adder.U$$681/X sky130_fd_sc_hd__a21o_1
XTAP_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_36_1 dadda_fa_3_36_1/A dadda_fa_3_36_1/B dadda_fa_3_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_0/CIN dadda_fa_4_36_2/A sky130_fd_sc_hd__fa_1
XU$$520 U$$520/A U$$528/B VGND VGND VPWR VPWR U$$520/X sky130_fd_sc_hd__xor2_1
XTAP_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$692 final_adder.U$$708/B final_adder.U$$692/B VGND VGND VPWR VPWR
+ final_adder.U$$772/A sky130_fd_sc_hd__and2_1
XTAP_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$531 U$$940/B1 U$$537/A2 U$$807/A1 U$$537/B2 VGND VGND VPWR VPWR U$$532/A sky130_fd_sc_hd__a22o_1
XFILLER_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_13_0 dadda_fa_6_13_0/A dadda_fa_6_13_0/B dadda_fa_6_13_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_14_0/B dadda_fa_7_13_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$542 U$$542/A U$$546/B VGND VGND VPWR VPWR U$$542/X sky130_fd_sc_hd__xor2_1
XTAP_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$553 U$$551/B U$$548/A U$$549/A U$$548/Y VGND VGND VPWR VPWR U$$553/X sky130_fd_sc_hd__a22o_4
XU$$564 U$$975/A1 U$$578/A2 U$$703/A1 U$$578/B2 VGND VGND VPWR VPWR U$$565/A sky130_fd_sc_hd__a22o_1
XTAP_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_29_0 U$$1528/X U$$1661/X U$$1794/X VGND VGND VPWR VPWR dadda_fa_4_30_0/B
+ dadda_fa_4_29_1/CIN sky130_fd_sc_hd__fa_1
XU$$575 U$$575/A U$$607/B VGND VGND VPWR VPWR U$$575/X sky130_fd_sc_hd__xor2_1
XFILLER_204_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$586 U$$721/B1 U$$606/A2 U$$40/A1 U$$606/B2 VGND VGND VPWR VPWR U$$587/A sky130_fd_sc_hd__a22o_1
XFILLER_16_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$597 U$$597/A U$$617/B VGND VGND VPWR VPWR U$$597/X sky130_fd_sc_hd__xor2_1
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_95_5 input251/X dadda_fa_2_95_5/B dadda_fa_2_95_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_96_2/A dadda_fa_4_95_0/A sky130_fd_sc_hd__fa_2
Xrepeater1420 U$$1870/B VGND VGND VPWR VPWR U$$1820/B sky130_fd_sc_hd__buf_6
XFILLER_67_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1431 input18/X VGND VGND VPWR VPWR U$$1779/B sky130_fd_sc_hd__buf_6
XFILLER_67_1023 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1442 U$$1592/B VGND VGND VPWR VPWR U$$1558/B sky130_fd_sc_hd__buf_8
Xrepeater1453 U$$1499/B VGND VGND VPWR VPWR U$$1501/B sky130_fd_sc_hd__buf_12
Xrepeater1464 input128/X VGND VGND VPWR VPWR U$$3451/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_88_4 dadda_fa_2_88_4/A dadda_fa_2_88_4/B dadda_fa_2_88_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_1/CIN dadda_fa_3_88_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_193_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1475 U$$3447/A1 VGND VGND VPWR VPWR U$$981/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1486 U$$431/A1 VGND VGND VPWR VPWR U$$20/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_207_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1497 U$$3555/B1 VGND VGND VPWR VPWR U$$3281/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_154_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_2_25_1 U$$456/X U$$589/X VGND VGND VPWR VPWR dadda_fa_3_26_3/A dadda_fa_4_25_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_31_0 U$$69/X U$$202/X U$$335/X VGND VGND VPWR VPWR dadda_fa_3_32_0/CIN
+ dadda_fa_3_31_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_51_923 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1270 U$$1270/A U$$1270/B VGND VGND VPWR VPWR U$$1270/X sky130_fd_sc_hd__xor2_1
XU$$1281 U$$733/A1 U$$1289/A2 U$$598/A1 U$$1281/B2 VGND VGND VPWR VPWR U$$1282/A sky130_fd_sc_hd__a22o_1
XFILLER_195_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1292 U$$1292/A U$$1330/B VGND VGND VPWR VPWR U$$1292/X sky130_fd_sc_hd__xor2_1
XFILLER_188_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_118_0 dadda_fa_5_118_0/A dadda_fa_5_118_0/B dadda_fa_5_118_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_119_0/A dadda_fa_6_118_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_3 U$$2567/X U$$2700/X U$$2833/X VGND VGND VPWR VPWR dadda_fa_2_84_2/CIN
+ dadda_fa_2_83_5/A sky130_fd_sc_hd__fa_1
XFILLER_46_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_60_2 dadda_fa_4_60_2/A dadda_fa_4_60_2/B dadda_fa_4_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_61_0/CIN dadda_fa_5_60_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_76_2 U$$2287/X U$$2420/X U$$2553/X VGND VGND VPWR VPWR dadda_fa_2_77_1/A
+ dadda_fa_2_76_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_53_1 dadda_fa_4_53_1/A dadda_fa_4_53_1/B dadda_fa_4_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/B dadda_fa_5_53_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_69_1 U$$2805/X U$$2938/X U$$3071/X VGND VGND VPWR VPWR dadda_fa_2_70_0/CIN
+ dadda_fa_2_69_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_30_0 dadda_fa_7_30_0/A dadda_fa_7_30_0/B dadda_fa_7_30_0/CIN VGND VGND
+ VPWR VPWR _327_/D _198_/D sky130_fd_sc_hd__fa_2
XFILLER_85_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_46_0 dadda_fa_4_46_0/A dadda_fa_4_46_0/B dadda_fa_4_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/A dadda_fa_5_46_1/A sky130_fd_sc_hd__fa_1
XFILLER_58_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_886 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _199_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_226 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_248 _292_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_259 U$$2302/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_361_ _362_/CLK _361_/D VGND VGND VPWR VPWR _361_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ _420_/CLK _292_/D VGND VGND VPWR VPWR _292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_98_3 dadda_fa_3_98_3/A dadda_fa_3_98_3/B dadda_fa_3_98_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_99_1/B dadda_fa_4_98_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_72_3 U$$1747/X U$$1880/X VGND VGND VPWR VPWR dadda_fa_1_73_8/A dadda_fa_2_72_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_5_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_71_1 U$$947/X U$$1080/X U$$1213/X VGND VGND VPWR VPWR dadda_fa_1_72_7/A
+ dadda_fa_1_71_8/B sky130_fd_sc_hd__fa_1
XFILLER_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_64_0 U$$135/X U$$268/X U$$401/X VGND VGND VPWR VPWR dadda_fa_1_65_5/B
+ dadda_fa_1_64_7/B sky130_fd_sc_hd__fa_1
XTAP_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$350 U$$76/A1 U$$350/A2 U$$78/A1 U$$350/B2 VGND VGND VPWR VPWR U$$351/A sky130_fd_sc_hd__a22o_1
XFILLER_205_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$361 U$$361/A U$$397/B VGND VGND VPWR VPWR U$$361/X sky130_fd_sc_hd__xor2_1
XFILLER_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$372 U$$920/A1 U$$378/A2 U$$920/B1 U$$378/B2 VGND VGND VPWR VPWR U$$373/A sky130_fd_sc_hd__a22o_1
XU$$383 U$$383/A U$$395/B VGND VGND VPWR VPWR U$$383/X sky130_fd_sc_hd__xor2_1
XFILLER_33_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$394 U$$942/A1 U$$394/A2 U$$944/A1 U$$394/B2 VGND VGND VPWR VPWR U$$395/A sky130_fd_sc_hd__a22o_1
XFILLER_60_775 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_93_2 U$$3651/X U$$3784/X U$$3917/X VGND VGND VPWR VPWR dadda_fa_3_94_1/A
+ dadda_fa_3_93_3/A sky130_fd_sc_hd__fa_1
XFILLER_161_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1250 U$$4080/B VGND VGND VPWR VPWR U$$4078/B sky130_fd_sc_hd__buf_6
Xdadda_fa_5_70_1 dadda_fa_5_70_1/A dadda_fa_5_70_1/B dadda_fa_5_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_71_0/B dadda_fa_7_70_0/A sky130_fd_sc_hd__fa_1
XFILLER_126_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_86_1 U$$4169/X U$$4302/X U$$4435/X VGND VGND VPWR VPWR dadda_fa_3_87_0/CIN
+ dadda_fa_3_86_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater1261 U$$3971/B VGND VGND VPWR VPWR U$$3972/A sky130_fd_sc_hd__buf_8
XFILLER_113_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1272 U$$3834/B VGND VGND VPWR VPWR U$$3814/B sky130_fd_sc_hd__buf_6
Xrepeater1283 U$$959/A VGND VGND VPWR VPWR U$$958/A sky130_fd_sc_hd__buf_12
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_63_0 dadda_fa_5_63_0/A dadda_fa_5_63_0/B dadda_fa_5_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_64_0/A dadda_fa_6_63_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1294 U$$3480/B VGND VGND VPWR VPWR U$$3454/B sky130_fd_sc_hd__buf_8
XFILLER_114_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_79_0 dadda_fa_2_79_0/A dadda_fa_2_79_0/B dadda_fa_2_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_0/B dadda_fa_3_79_2/B sky130_fd_sc_hd__fa_1
XFILLER_59_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1110 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_62_8 dadda_fa_1_62_8/A dadda_fa_1_62_8/B dadda_fa_1_62_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_63_3/A dadda_fa_3_62_0/A sky130_fd_sc_hd__fa_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_55_7 U$$3575/X U$$3708/X input207/X VGND VGND VPWR VPWR dadda_fa_2_56_2/CIN
+ dadda_fa_2_55_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_48_6 U$$2497/X U$$2630/X U$$2763/X VGND VGND VPWR VPWR dadda_fa_2_49_3/A
+ dadda_fa_2_48_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_167_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_56 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_78_0 dadda_fa_7_78_0/A dadda_fa_7_78_0/B dadda_fa_7_78_0/CIN VGND VGND
+ VPWR VPWR _375_/D _246_/D sky130_fd_sc_hd__fa_1
XFILLER_192_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_81_0 U$$1232/Y U$$1366/X U$$1499/X VGND VGND VPWR VPWR dadda_fa_2_82_1/A
+ dadda_fa_2_81_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_144_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4109 U$$4109/A VGND VGND VPWR VPWR U$$4109/Y sky130_fd_sc_hd__inv_1
XFILLER_120_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3408 U$$3545/A1 U$$3422/A2 U$$3684/A1 U$$3422/B2 VGND VGND VPWR VPWR U$$3409/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3419 U$$3419/A U$$3424/A VGND VGND VPWR VPWR U$$3419/X sky130_fd_sc_hd__xor2_1
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2707 U$$2842/B1 U$$2607/X U$$2709/A1 U$$2608/X VGND VGND VPWR VPWR U$$2708/A sky130_fd_sc_hd__a22o_1
XFILLER_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2718 U$$2718/A U$$2739/A VGND VGND VPWR VPWR U$$2718/X sky130_fd_sc_hd__xor2_1
XFILLER_46_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2729 U$$3414/A1 U$$2735/A2 U$$3414/B1 U$$2735/B2 VGND VGND VPWR VPWR U$$2730/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_413_ _414_/CLK _413_/D VGND VGND VPWR VPWR _413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_344_ _351_/CLK _344_/D VGND VGND VPWR VPWR _344_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_499 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_275_ _407_/CLK _275_/D VGND VGND VPWR VPWR _275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_80_0 dadda_fa_6_80_0/A dadda_fa_6_80_0/B dadda_fa_6_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_81_0/B dadda_fa_7_80_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_96_0 dadda_fa_3_96_0/A dadda_fa_3_96_0/B dadda_fa_3_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_0/B dadda_fa_4_96_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater906 U$$2691/A1 VGND VGND VPWR VPWR U$$2415/B1 sky130_fd_sc_hd__buf_6
Xrepeater917 input98/X VGND VGND VPWR VPWR U$$3300/B1 sky130_fd_sc_hd__buf_6
XFILLER_209_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater928 U$$2550/A1 VGND VGND VPWR VPWR U$$630/B1 sky130_fd_sc_hd__buf_4
Xrepeater939 U$$3368/B1 VGND VGND VPWR VPWR U$$2409/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_58_5 dadda_fa_2_58_5/A dadda_fa_2_58_5/B dadda_fa_2_58_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_2/A dadda_fa_4_58_0/A sky130_fd_sc_hd__fa_2
XFILLER_76_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3920 U$$4055/B1 U$$3926/A2 U$$4333/A1 U$$3926/B2 VGND VGND VPWR VPWR U$$3921/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3931 U$$3931/A U$$3947/B VGND VGND VPWR VPWR U$$3931/X sky130_fd_sc_hd__xor2_1
XTAP_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3942 U$$4077/B1 U$$3946/A2 U$$3944/A1 U$$3946/B2 VGND VGND VPWR VPWR U$$3943/A
+ sky130_fd_sc_hd__a22o_1
XU$$3953 U$$3953/A U$$3972/A VGND VGND VPWR VPWR U$$3953/X sky130_fd_sc_hd__xor2_1
XTAP_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3964 U$$4512/A1 U$$3968/A2 U$$4240/A1 U$$3968/B2 VGND VGND VPWR VPWR U$$3965/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_840 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3975 U$$4109/A VGND VGND VPWR VPWR U$$3975/Y sky130_fd_sc_hd__inv_1
XFILLER_18_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3986 U$$3986/A U$$4044/B VGND VGND VPWR VPWR U$$3986/X sky130_fd_sc_hd__xor2_1
XU$$3997 U$$4408/A1 U$$4035/A2 U$$4273/A1 U$$4035/B2 VGND VGND VPWR VPWR U$$3998/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$180 U$$180/A U$$212/B VGND VGND VPWR VPWR U$$180/X sky130_fd_sc_hd__xor2_1
XU$$191 U$$328/A1 U$$217/A2 U$$328/B1 U$$217/B2 VGND VGND VPWR VPWR U$$192/A sky130_fd_sc_hd__a22o_1
XFILLER_21_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput266 output266/A VGND VGND VPWR VPWR o[108] sky130_fd_sc_hd__buf_2
Xrepeater1080 U$$4162/A1 VGND VGND VPWR VPWR U$$4297/B1 sky130_fd_sc_hd__clkbuf_8
Xoutput277 output277/A VGND VGND VPWR VPWR o[118] sky130_fd_sc_hd__buf_2
XFILLER_134_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1091 U$$4293/B1 VGND VGND VPWR VPWR U$$3473/A1 sky130_fd_sc_hd__buf_6
Xoutput288 output288/A VGND VGND VPWR VPWR o[12] sky130_fd_sc_hd__buf_2
XFILLER_88_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput299 output299/A VGND VGND VPWR VPWR o[22] sky130_fd_sc_hd__buf_2
XFILLER_82_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_60_5 U$$3984/X U$$4117/X U$$4145/B VGND VGND VPWR VPWR dadda_fa_2_61_2/A
+ dadda_fa_2_60_5/A sky130_fd_sc_hd__fa_1
XFILLER_101_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_4 U$$1975/X U$$2108/X U$$2241/X VGND VGND VPWR VPWR dadda_fa_2_54_1/CIN
+ dadda_fa_2_53_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_46_3 U$$1296/X U$$1429/X U$$1562/X VGND VGND VPWR VPWR dadda_fa_2_47_2/CIN
+ dadda_fa_2_46_5/A sky130_fd_sc_hd__fa_1
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_23_2 dadda_fa_4_23_2/A dadda_fa_4_23_2/B dadda_fa_4_23_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_24_0/CIN dadda_fa_5_23_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_16_1 U$$1103/X U$$1139/B input164/X VGND VGND VPWR VPWR dadda_fa_5_17_0/B
+ dadda_fa_5_16_1/B sky130_fd_sc_hd__fa_1
XFILLER_180_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_747 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1107 final_adder.U$$172/B final_adder.U$$943/X VGND VGND VPWR VPWR
+ output366/A sky130_fd_sc_hd__xor2_1
XFILLER_104_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1118 final_adder.U$$160/A final_adder.U$$869/X VGND VGND VPWR VPWR
+ output378/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1129 final_adder.U$$150/B final_adder.U$$921/X VGND VGND VPWR VPWR
+ output263/A sky130_fd_sc_hd__xor2_1
XFILLER_20_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1048 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1062 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3205 U$$4162/B1 U$$3207/A2 U$$4440/A1 U$$3207/B2 VGND VGND VPWR VPWR U$$3206/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3216 U$$3216/A U$$3228/B VGND VGND VPWR VPWR U$$3216/X sky130_fd_sc_hd__xor2_1
XFILLER_171_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3227 U$$3775/A1 U$$3229/A2 U$$3775/B1 U$$3227/B2 VGND VGND VPWR VPWR U$$3228/A
+ sky130_fd_sc_hd__a22o_1
XU$$3238 U$$3238/A U$$3242/B VGND VGND VPWR VPWR U$$3238/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2504 U$$312/A1 U$$2596/A2 U$$38/B1 U$$2596/B2 VGND VGND VPWR VPWR U$$2505/A sky130_fd_sc_hd__a22o_1
XU$$3249 U$$4480/B1 U$$3285/A2 U$$4484/A1 U$$3285/B2 VGND VGND VPWR VPWR U$$3250/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2515 U$$2515/A U$$2601/B VGND VGND VPWR VPWR U$$2515/X sky130_fd_sc_hd__xor2_1
XU$$2526 U$$2661/B1 U$$2558/A2 U$$62/A1 U$$2558/B2 VGND VGND VPWR VPWR U$$2527/A sky130_fd_sc_hd__a22o_1
XFILLER_74_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2537 U$$2537/A U$$2543/B VGND VGND VPWR VPWR U$$2537/X sky130_fd_sc_hd__xor2_1
XFILLER_34_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2548 U$$2683/B1 U$$2600/A2 U$$2550/A1 U$$2600/B2 VGND VGND VPWR VPWR U$$2549/A
+ sky130_fd_sc_hd__a22o_1
XU$$1803 U$$981/A1 U$$1839/A2 U$$709/A1 U$$1839/B2 VGND VGND VPWR VPWR U$$1804/A sky130_fd_sc_hd__a22o_1
XU$$1814 U$$1814/A U$$1820/B VGND VGND VPWR VPWR U$$1814/X sky130_fd_sc_hd__xor2_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2559 U$$2559/A U$$2569/B VGND VGND VPWR VPWR U$$2559/X sky130_fd_sc_hd__xor2_1
XFILLER_203_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1825 U$$3058/A1 U$$1877/A2 U$$3606/B1 U$$1877/B2 VGND VGND VPWR VPWR U$$1826/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1836 U$$1836/A U$$1840/B VGND VGND VPWR VPWR U$$1836/X sky130_fd_sc_hd__xor2_1
XFILLER_187_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1847 U$$1984/A1 U$$1879/A2 U$$2123/A1 U$$1879/B2 VGND VGND VPWR VPWR U$$1848/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1858 U$$1858/A U$$1870/B VGND VGND VPWR VPWR U$$1858/X sky130_fd_sc_hd__xor2_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1869 U$$2691/A1 U$$1869/A2 U$$2282/A1 U$$1869/B2 VGND VGND VPWR VPWR U$$1870/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_327_ _327_/CLK _327_/D VGND VGND VPWR VPWR _327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_258_ _387_/CLK _258_/D VGND VGND VPWR VPWR _258_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_190_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_189_ _327_/CLK _189_/D VGND VGND VPWR VPWR _189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_70_4 dadda_fa_2_70_4/A dadda_fa_2_70_4/B dadda_fa_2_70_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_1/CIN dadda_fa_3_70_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_63_3 dadda_fa_2_63_3/A dadda_fa_2_63_3/B dadda_fa_2_63_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/B dadda_fa_3_63_3/B sky130_fd_sc_hd__fa_1
Xrepeater703 U$$3874/B2 VGND VGND VPWR VPWR U$$3902/B2 sky130_fd_sc_hd__buf_6
XFILLER_85_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater714 U$$3777/B2 VGND VGND VPWR VPWR U$$3833/B2 sky130_fd_sc_hd__buf_6
XFILLER_111_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater725 U$$3567/X VGND VGND VPWR VPWR U$$3636/B2 sky130_fd_sc_hd__buf_4
XFILLER_111_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_56_2 dadda_fa_2_56_2/A dadda_fa_2_56_2/B dadda_fa_2_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/A dadda_fa_3_56_3/A sky130_fd_sc_hd__fa_1
Xrepeater736 U$$3378/B2 VGND VGND VPWR VPWR U$$3346/B2 sky130_fd_sc_hd__buf_6
XFILLER_84_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater747 U$$3285/B2 VGND VGND VPWR VPWR U$$3277/B2 sky130_fd_sc_hd__buf_4
XFILLER_38_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater758 U$$2985/B2 VGND VGND VPWR VPWR U$$2995/B2 sky130_fd_sc_hd__buf_4
XU$$4440 U$$4440/A1 U$$4388/X U$$4440/B1 U$$4389/X VGND VGND VPWR VPWR U$$4441/A sky130_fd_sc_hd__a22o_1
XFILLER_93_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_33_1 dadda_fa_5_33_1/A dadda_fa_5_33_1/B dadda_fa_5_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_34_0/B dadda_fa_7_33_0/A sky130_fd_sc_hd__fa_1
Xrepeater769 U$$366/B2 VGND VGND VPWR VPWR U$$340/B2 sky130_fd_sc_hd__buf_4
XU$$4451 U$$4451/A U$$4451/B VGND VGND VPWR VPWR U$$4451/X sky130_fd_sc_hd__xor2_1
XFILLER_42_1187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4462 input93/X U$$4388/X U$$4464/A1 U$$4476/B2 VGND VGND VPWR VPWR U$$4463/A sky130_fd_sc_hd__a22o_1
XFILLER_37_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_49_1 dadda_fa_2_49_1/A dadda_fa_2_49_1/B dadda_fa_2_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_0/CIN dadda_fa_3_49_2/CIN sky130_fd_sc_hd__fa_1
XU$$4473 U$$4473/A U$$4473/B VGND VGND VPWR VPWR U$$4473/X sky130_fd_sc_hd__xor2_1
XU$$4484 U$$4484/A1 U$$4388/X U$$4484/B1 U$$4486/B2 VGND VGND VPWR VPWR U$$4485/A
+ sky130_fd_sc_hd__a22o_1
XU$$3750 U$$3750/A U$$3794/B VGND VGND VPWR VPWR U$$3750/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_26_0 dadda_fa_5_26_0/A dadda_fa_5_26_0/B dadda_fa_5_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_27_0/A dadda_fa_6_26_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_77_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4495 U$$4495/A U$$4495/B VGND VGND VPWR VPWR U$$4495/X sky130_fd_sc_hd__xor2_1
XFILLER_25_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3761 U$$3761/A1 U$$3703/X U$$4311/A1 U$$3704/X VGND VGND VPWR VPWR U$$3762/A sky130_fd_sc_hd__a22o_1
XU$$3772 U$$3772/A U$$3774/B VGND VGND VPWR VPWR U$$3772/X sky130_fd_sc_hd__xor2_1
XFILLER_53_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3783 U$$4466/B1 U$$3813/A2 U$$4468/B1 U$$3813/B2 VGND VGND VPWR VPWR U$$3784/A
+ sky130_fd_sc_hd__a22o_1
XU$$3794 U$$3794/A U$$3794/B VGND VGND VPWR VPWR U$$3794/X sky130_fd_sc_hd__xor2_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_100_0 dadda_fa_5_100_0/A dadda_fa_5_100_0/B dadda_fa_5_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_101_0/A dadda_fa_6_100_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_146_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_992 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_51_1 U$$508/X U$$641/X U$$774/X VGND VGND VPWR VPWR dadda_fa_2_52_0/CIN
+ dadda_fa_2_51_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_141_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$905 U$$905/A U$$951/B VGND VGND VPWR VPWR U$$905/X sky130_fd_sc_hd__xor2_1
XFILLER_55_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$916 U$$916/A1 U$$918/A2 U$$916/B1 U$$918/B2 VGND VGND VPWR VPWR U$$917/A sky130_fd_sc_hd__a22o_1
XFILLER_84_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_44_0 U$$95/X U$$228/X U$$361/X VGND VGND VPWR VPWR dadda_fa_2_45_2/B dadda_fa_2_44_4/B
+ sky130_fd_sc_hd__fa_1
XU$$927 U$$927/A U$$945/B VGND VGND VPWR VPWR U$$927/X sky130_fd_sc_hd__xor2_1
XFILLER_56_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$938 U$$938/A1 U$$938/A2 U$$940/A1 U$$938/B2 VGND VGND VPWR VPWR U$$939/A sky130_fd_sc_hd__a22o_1
XFILLER_16_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$949 U$$949/A U$$958/A VGND VGND VPWR VPWR U$$949/X sky130_fd_sc_hd__xor2_1
XFILLER_189_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_634 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_892 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1069 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_80_3 dadda_fa_3_80_3/A dadda_fa_3_80_3/B dadda_fa_3_80_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_1/B dadda_fa_4_80_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_65_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_73_2 dadda_fa_3_73_2/A dadda_fa_3_73_2/B dadda_fa_3_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_1/A dadda_fa_4_73_2/B sky130_fd_sc_hd__fa_1
XFILLER_191_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_66_1 dadda_fa_3_66_1/A dadda_fa_3_66_1/B dadda_fa_3_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_0/CIN dadda_fa_4_66_2/A sky130_fd_sc_hd__fa_1
XU$$4415_1784 VGND VGND VPWR VPWR U$$4415_1784/HI U$$4415/B sky130_fd_sc_hd__conb_1
XFILLER_26_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_43_0 dadda_fa_6_43_0/A dadda_fa_6_43_0/B dadda_fa_6_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_44_0/B dadda_fa_7_43_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_59_0 dadda_fa_3_59_0/A dadda_fa_3_59_0/B dadda_fa_3_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_0/B dadda_fa_4_59_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3002 U$$3002/A U$$3013/A VGND VGND VPWR VPWR U$$3002/X sky130_fd_sc_hd__xor2_1
XFILLER_208_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3013 U$$3013/A VGND VGND VPWR VPWR U$$3013/Y sky130_fd_sc_hd__inv_1
XFILLER_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3024 U$$3159/B1 U$$3060/A2 U$$4396/A1 U$$3060/B2 VGND VGND VPWR VPWR U$$3025/A
+ sky130_fd_sc_hd__a22o_1
XU$$3035 U$$3035/A U$$3083/B VGND VGND VPWR VPWR U$$3035/X sky130_fd_sc_hd__xor2_1
XU$$3046 input68/X U$$3124/A2 U$$32/B1 U$$3124/B2 VGND VGND VPWR VPWR U$$3047/A sky130_fd_sc_hd__a22o_1
XFILLER_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2301 U$$2301/A input27/X VGND VGND VPWR VPWR U$$2301/X sky130_fd_sc_hd__xor2_1
XFILLER_74_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3057 U$$3057/A U$$3075/B VGND VGND VPWR VPWR U$$3057/X sky130_fd_sc_hd__xor2_1
XU$$2312 U$$2312/A1 U$$2196/X U$$2312/B1 U$$2197/X VGND VGND VPWR VPWR U$$2313/A sky130_fd_sc_hd__a22o_1
XFILLER_75_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_102_2 dadda_fa_4_102_2/A dadda_fa_4_102_2/B dadda_fa_4_102_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_103_0/CIN dadda_fa_5_102_1/CIN sky130_fd_sc_hd__fa_1
XU$$2323 U$$2323/A U$$2328/A VGND VGND VPWR VPWR U$$2323/X sky130_fd_sc_hd__xor2_1
XFILLER_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3068 U$$4162/B1 U$$3098/A2 U$$3344/A1 U$$3098/B2 VGND VGND VPWR VPWR U$$3069/A
+ sky130_fd_sc_hd__a22o_1
XU$$2334 U$$2332/B input27/X input28/X U$$2329/Y VGND VGND VPWR VPWR U$$2334/X sky130_fd_sc_hd__a22o_4
XFILLER_90_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1600 U$$1600/A U$$1608/B VGND VGND VPWR VPWR U$$1600/X sky130_fd_sc_hd__xor2_1
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3079 U$$3079/A U$$3083/B VGND VGND VPWR VPWR U$$3079/X sky130_fd_sc_hd__xor2_1
XU$$2345 U$$2754/B1 U$$2359/A2 U$$2621/A1 U$$2359/B2 VGND VGND VPWR VPWR U$$2346/A
+ sky130_fd_sc_hd__a22o_1
XU$$2356 U$$2356/A U$$2360/B VGND VGND VPWR VPWR U$$2356/X sky130_fd_sc_hd__xor2_1
XU$$1611 U$$2568/B1 U$$1635/A2 U$$2159/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1612/A
+ sky130_fd_sc_hd__a22o_1
XU$$2367 U$$312/A1 U$$2463/A2 U$$40/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2368/A sky130_fd_sc_hd__a22o_1
XFILLER_37_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1622 U$$1622/A U$$1628/B VGND VGND VPWR VPWR U$$1622/X sky130_fd_sc_hd__xor2_1
XU$$2378 U$$2378/A U$$2380/B VGND VGND VPWR VPWR U$$2378/X sky130_fd_sc_hd__xor2_1
XFILLER_22_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1633 U$$948/A1 U$$1637/A2 U$$950/A1 U$$1637/B2 VGND VGND VPWR VPWR U$$1634/A sky130_fd_sc_hd__a22o_1
XFILLER_76_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1644 U$$1644/A VGND VGND VPWR VPWR U$$1644/Y sky130_fd_sc_hd__inv_1
XU$$2389 U$$882/A1 U$$2403/A2 U$$2391/A1 U$$2403/B2 VGND VGND VPWR VPWR U$$2390/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1655 U$$1655/A U$$1689/B VGND VGND VPWR VPWR U$$1655/X sky130_fd_sc_hd__xor2_1
XFILLER_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1666 U$$1666/A1 U$$1696/A2 U$$1666/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1667/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1677 U$$1677/A U$$1679/B VGND VGND VPWR VPWR U$$1677/X sky130_fd_sc_hd__xor2_1
XFILLER_203_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1688 U$$727/B1 U$$1688/A2 U$$594/A1 U$$1688/B2 VGND VGND VPWR VPWR U$$1689/A sky130_fd_sc_hd__a22o_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1699 U$$1699/A U$$1751/B VGND VGND VPWR VPWR U$$1699/X sky130_fd_sc_hd__xor2_1
XFILLER_175_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_116_0 dadda_fa_7_116_0/A dadda_fa_7_116_0/B dadda_fa_7_116_0/CIN VGND
+ VGND VPWR VPWR _413_/D _284_/D sky130_fd_sc_hd__fa_1
XFILLER_204_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_61_0 dadda_fa_2_61_0/A dadda_fa_2_61_0/B dadda_fa_2_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_0/B dadda_fa_3_61_2/B sky130_fd_sc_hd__fa_1
Xrepeater500 U$$3241/A2 VGND VGND VPWR VPWR U$$3207/A2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$307 final_adder.U$$306/B final_adder.U$$181/X final_adder.U$$179/X
+ VGND VGND VPWR VPWR final_adder.U$$307/X sky130_fd_sc_hd__a21o_1
Xrepeater511 U$$2985/A2 VGND VGND VPWR VPWR U$$2995/A2 sky130_fd_sc_hd__buf_4
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$318 final_adder.U$$320/B final_adder.U$$318/B VGND VGND VPWR VPWR
+ final_adder.U$$444/B sky130_fd_sc_hd__and2_1
Xrepeater522 U$$366/A2 VGND VGND VPWR VPWR U$$340/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$329 final_adder.U$$328/B final_adder.U$$203/X final_adder.U$$201/X
+ VGND VGND VPWR VPWR final_adder.U$$329/X sky130_fd_sc_hd__a21o_1
Xrepeater533 U$$2828/A2 VGND VGND VPWR VPWR U$$2874/A2 sky130_fd_sc_hd__buf_6
Xrepeater544 U$$2600/A2 VGND VGND VPWR VPWR U$$2596/A2 sky130_fd_sc_hd__clkbuf_8
Xrepeater555 U$$2449/A2 VGND VGND VPWR VPWR U$$2435/A2 sky130_fd_sc_hd__buf_6
XFILLER_38_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater566 U$$2196/X VGND VGND VPWR VPWR U$$2302/A2 sky130_fd_sc_hd__buf_6
Xrepeater577 U$$2016/A2 VGND VGND VPWR VPWR U$$1990/A2 sky130_fd_sc_hd__buf_8
Xrepeater588 U$$1913/A2 VGND VGND VPWR VPWR U$$1879/A2 sky130_fd_sc_hd__buf_4
XU$$4270 U$$4270/A U$$4278/B VGND VGND VPWR VPWR U$$4270/X sky130_fd_sc_hd__xor2_1
XU$$4281 input69/X U$$4327/A2 input70/X U$$4327/B2 VGND VGND VPWR VPWR U$$4282/A sky130_fd_sc_hd__a22o_1
Xrepeater599 U$$1648/X VGND VGND VPWR VPWR U$$1770/A2 sky130_fd_sc_hd__buf_6
XFILLER_53_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4292 U$$4292/A U$$4294/B VGND VGND VPWR VPWR U$$4292/X sky130_fd_sc_hd__xor2_1
XFILLER_77_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3580 input120/X U$$3612/A2 U$$4404/A1 U$$3612/B2 VGND VGND VPWR VPWR U$$3581/A
+ sky130_fd_sc_hd__a22o_1
XU$$3591 U$$3591/A U$$3613/B VGND VGND VPWR VPWR U$$3591/X sky130_fd_sc_hd__xor2_1
XFILLER_41_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2890 U$$2890/A U$$2922/B VGND VGND VPWR VPWR U$$2890/X sky130_fd_sc_hd__xor2_1
XFILLER_178_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_90_2 dadda_fa_4_90_2/A dadda_fa_4_90_2/B dadda_fa_4_90_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_91_0/CIN dadda_fa_5_90_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_179_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_83_1 dadda_fa_4_83_1/A dadda_fa_4_83_1/B dadda_fa_4_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/B dadda_fa_5_83_1/B sky130_fd_sc_hd__fa_1
XFILLER_134_444 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_60_0 dadda_fa_7_60_0/A dadda_fa_7_60_0/B dadda_fa_7_60_0/CIN VGND VGND
+ VPWR VPWR _357_/D _228_/D sky130_fd_sc_hd__fa_1
XFILLER_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_76_0 dadda_fa_4_76_0/A dadda_fa_4_76_0/B dadda_fa_4_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/A dadda_fa_5_76_1/A sky130_fd_sc_hd__fa_1
XFILLER_161_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$841 final_adder.U$$744/X final_adder.U$$809/X final_adder.U$$745/X
+ VGND VGND VPWR VPWR final_adder.U$$841/X sky130_fd_sc_hd__a21o_2
XTAP_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$863 final_adder.U$$766/X final_adder.U$$831/X final_adder.U$$767/X
+ VGND VGND VPWR VPWR final_adder.U$$863/X sky130_fd_sc_hd__a21o_2
XTAP_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$702 U$$702/A U$$712/B VGND VGND VPWR VPWR U$$702/X sky130_fd_sc_hd__xor2_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$713 U$$850/A1 U$$739/A2 U$$850/B1 U$$739/B2 VGND VGND VPWR VPWR U$$714/A sky130_fd_sc_hd__a22o_1
XFILLER_1_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$885 final_adder.U$$788/X final_adder.U$$621/X final_adder.U$$789/X
+ VGND VGND VPWR VPWR final_adder.U$$885/X sky130_fd_sc_hd__a21o_1
XU$$724 U$$724/A U$$750/B VGND VGND VPWR VPWR U$$724/X sky130_fd_sc_hd__xor2_1
XFILLER_90_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$735 U$$48/B1 U$$749/A2 U$$52/A1 U$$749/B2 VGND VGND VPWR VPWR U$$736/A sky130_fd_sc_hd__a22o_1
XU$$746 U$$746/A U$$750/B VGND VGND VPWR VPWR U$$746/X sky130_fd_sc_hd__xor2_1
XU$$757 U$$757/A1 U$$759/A2 U$$896/A1 U$$759/B2 VGND VGND VPWR VPWR U$$758/A sky130_fd_sc_hd__a22o_1
XFILLER_44_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$768 U$$768/A U$$770/B VGND VGND VPWR VPWR U$$768/X sky130_fd_sc_hd__xor2_1
XU$$779 U$$914/B1 U$$783/A2 U$$918/A1 U$$783/B2 VGND VGND VPWR VPWR U$$780/A sky130_fd_sc_hd__a22o_1
XFILLER_72_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_639 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4445_1799 VGND VGND VPWR VPWR U$$4445_1799/HI U$$4445/B sky130_fd_sc_hd__conb_1
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1602 input112/X VGND VGND VPWR VPWR U$$4496/A1 sky130_fd_sc_hd__buf_6
XANTENNA_7 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1613 U$$2848/A1 VGND VGND VPWR VPWR U$$2026/A1 sky130_fd_sc_hd__buf_4
Xrepeater1624 U$$1316/B VGND VGND VPWR VPWR U$$1272/B sky130_fd_sc_hd__buf_6
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1635 U$$3852/A1 VGND VGND VPWR VPWR U$$3987/B1 sky130_fd_sc_hd__buf_4
XFILLER_125_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1646 U$$3801/B1 VGND VGND VPWR VPWR U$$652/A1 sky130_fd_sc_hd__buf_4
Xrepeater1657 U$$2292/B1 VGND VGND VPWR VPWR U$$924/A1 sky130_fd_sc_hd__buf_8
XFILLER_99_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1668 input105/X VGND VGND VPWR VPWR U$$4484/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1679 U$$4478/B1 VGND VGND VPWR VPWR U$$4343/A1 sky130_fd_sc_hd__buf_6
XFILLER_98_328 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1085 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_40_5 dadda_fa_2_40_5/A dadda_fa_2_40_5/B dadda_fa_2_40_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_41_2/A dadda_fa_4_40_0/A sky130_fd_sc_hd__fa_2
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_33_4 U$$1669/X U$$1802/X U$$1935/X VGND VGND VPWR VPWR dadda_fa_3_34_1/CIN
+ dadda_fa_3_33_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2120 U$$2120/A U$$2150/B VGND VGND VPWR VPWR U$$2120/X sky130_fd_sc_hd__xor2_1
XU$$2131 U$$896/B1 U$$2177/A2 U$$3366/A1 U$$2177/B2 VGND VGND VPWR VPWR U$$2132/A
+ sky130_fd_sc_hd__a22o_1
XU$$2142 U$$2142/A U$$2170/B VGND VGND VPWR VPWR U$$2142/X sky130_fd_sc_hd__xor2_1
XFILLER_90_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2153 U$$783/A1 U$$2189/A2 U$$920/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2154/A sky130_fd_sc_hd__a22o_1
XFILLER_90_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2164 U$$2164/A U$$2184/B VGND VGND VPWR VPWR U$$2164/X sky130_fd_sc_hd__xor2_1
XFILLER_179_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2175 U$$2312/A1 U$$2177/A2 U$$2312/B1 U$$2177/B2 VGND VGND VPWR VPWR U$$2176/A
+ sky130_fd_sc_hd__a22o_1
XU$$1430 U$$882/A1 U$$1434/A2 U$$2391/A1 U$$1434/B2 VGND VGND VPWR VPWR U$$1431/A
+ sky130_fd_sc_hd__a22o_1
XU$$2186 U$$2186/A U$$2191/A VGND VGND VPWR VPWR U$$2186/X sky130_fd_sc_hd__xor2_1
XU$$1441 U$$1441/A U$$1449/B VGND VGND VPWR VPWR U$$1441/X sky130_fd_sc_hd__xor2_1
XFILLER_16_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2197 U$$2195/B input25/X input26/X U$$2192/Y VGND VGND VPWR VPWR U$$2197/X sky130_fd_sc_hd__a22o_4
XU$$1452 U$$2683/B1 U$$1504/A2 U$$2550/A1 U$$1504/B2 VGND VGND VPWR VPWR U$$1453/A
+ sky130_fd_sc_hd__a22o_1
XU$$1463 U$$1463/A U$$1506/A VGND VGND VPWR VPWR U$$1463/X sky130_fd_sc_hd__xor2_1
XU$$1474 U$$2568/B1 U$$1374/X U$$2159/B1 U$$1375/X VGND VGND VPWR VPWR U$$1475/A sky130_fd_sc_hd__a22o_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1485 U$$1485/A U$$1501/B VGND VGND VPWR VPWR U$$1485/X sky130_fd_sc_hd__xor2_1
XFILLER_124_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1496 U$$4510/A1 U$$1502/A2 U$$2318/B1 U$$1502/B2 VGND VGND VPWR VPWR U$$1497/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_93_0 dadda_fa_5_93_0/A dadda_fa_5_93_0/B dadda_fa_5_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_94_0/A dadda_fa_6_93_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_204_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_78_6 U$$3621/X U$$3754/X U$$3887/X VGND VGND VPWR VPWR dadda_fa_2_79_2/B
+ dadda_fa_2_78_5/B sky130_fd_sc_hd__fa_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$104 _400_/Q _272_/Q VGND VGND VPWR VPWR final_adder.U$$921/B1 final_adder.U$$150/A
+ sky130_fd_sc_hd__ha_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$115 _411_/Q _283_/Q VGND VGND VPWR VPWR final_adder.U$$141/B1 final_adder.U$$140/B
+ sky130_fd_sc_hd__ha_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$126 _422_/Q _294_/Q VGND VGND VPWR VPWR final_adder.U$$899/B1 final_adder.U$$899/A1
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$137 final_adder.U$$136/B final_adder.U$$907/B1 final_adder.U$$137/B1
+ VGND VGND VPWR VPWR final_adder.U$$137/X sky130_fd_sc_hd__a21o_1
XFILLER_131_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$148 final_adder.U$$148/A final_adder.U$$148/B VGND VGND VPWR VPWR
+ final_adder.U$$276/B sky130_fd_sc_hd__and2_1
XTAP_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$159 final_adder.U$$158/B final_adder.U$$929/B1 final_adder.U$$159/B1
+ VGND VGND VPWR VPWR final_adder.U$$159/X sky130_fd_sc_hd__a21o_1
XFILLER_26_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater385 U$$1083/A2 VGND VGND VPWR VPWR U$$993/A2 sky130_fd_sc_hd__buf_4
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater396 U$$950/A2 VGND VGND VPWR VPWR U$$906/A2 sky130_fd_sc_hd__buf_4
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_102_1 U$$4467/X input132/X dadda_fa_3_102_1/CIN VGND VGND VPWR VPWR dadda_fa_4_103_0/CIN
+ dadda_fa_4_102_2/A sky130_fd_sc_hd__fa_2
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_274 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput100 b[41] VGND VGND VPWR VPWR input100/X sky130_fd_sc_hd__buf_6
Xinput111 b[51] VGND VGND VPWR VPWR input111/X sky130_fd_sc_hd__buf_6
XFILLER_153_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput122 b[61] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__buf_8
XFILLER_88_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_123_0 dadda_fa_6_123_0/A dadda_fa_6_123_0/B dadda_fa_6_123_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_124_0/B dadda_fa_7_123_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput133 c[103] VGND VGND VPWR VPWR input133/X sky130_fd_sc_hd__clkbuf_4
Xinput144 c[113] VGND VGND VPWR VPWR input144/X sky130_fd_sc_hd__buf_4
XFILLER_209_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput155 c[123] VGND VGND VPWR VPWR input155/X sky130_fd_sc_hd__buf_2
Xdadda_fa_0_66_4 U$$1735/X U$$1868/X U$$2001/X VGND VGND VPWR VPWR dadda_fa_1_67_6/CIN
+ dadda_fa_1_66_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 c[18] VGND VGND VPWR VPWR input166/X sky130_fd_sc_hd__clkbuf_4
XTAP_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput177 c[28] VGND VGND VPWR VPWR input177/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_43_3 dadda_fa_3_43_3/A dadda_fa_3_43_3/B dadda_fa_3_43_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_1/B dadda_fa_4_43_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 c[38] VGND VGND VPWR VPWR input188/X sky130_fd_sc_hd__clkbuf_2
XTAP_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput199 c[48] VGND VGND VPWR VPWR input199/X sky130_fd_sc_hd__clkbuf_2
Xfinal_adder.U$$660 final_adder.U$$676/B final_adder.U$$660/B VGND VGND VPWR VPWR
+ final_adder.U$$772/B sky130_fd_sc_hd__and2_1
XTAP_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$671 final_adder.U$$670/B final_adder.U$$567/X final_adder.U$$551/X
+ VGND VGND VPWR VPWR final_adder.U$$671/X sky130_fd_sc_hd__a21o_1
XTAP_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$510 U$$510/A U$$516/B VGND VGND VPWR VPWR U$$510/X sky130_fd_sc_hd__xor2_1
XFILLER_205_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$682 final_adder.U$$698/B final_adder.U$$682/B VGND VGND VPWR VPWR
+ final_adder.U$$794/B sky130_fd_sc_hd__and2_1
XTAP_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_36_2 dadda_fa_3_36_2/A dadda_fa_3_36_2/B dadda_fa_3_36_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_1/A dadda_fa_4_36_2/B sky130_fd_sc_hd__fa_1
XU$$521 U$$521/A1 U$$521/A2 U$$521/B1 U$$521/B2 VGND VGND VPWR VPWR U$$522/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$693 final_adder.U$$692/B final_adder.U$$589/X final_adder.U$$573/X
+ VGND VGND VPWR VPWR final_adder.U$$693/X sky130_fd_sc_hd__a21o_1
XTAP_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$532 U$$532/A U$$536/B VGND VGND VPWR VPWR U$$532/X sky130_fd_sc_hd__xor2_1
XFILLER_91_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$543 U$$678/B1 U$$415/X U$$817/B1 U$$416/X VGND VGND VPWR VPWR U$$544/A sky130_fd_sc_hd__a22o_1
XU$$554 U$$554/A1 U$$606/A2 U$$8/A1 U$$606/B2 VGND VGND VPWR VPWR U$$555/A sky130_fd_sc_hd__a22o_1
XTAP_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_29_1 U$$1927/X input178/X dadda_fa_3_29_1/CIN VGND VGND VPWR VPWR dadda_fa_4_30_0/CIN
+ dadda_fa_4_29_2/A sky130_fd_sc_hd__fa_1
XU$$565 U$$565/A U$$579/B VGND VGND VPWR VPWR U$$565/X sky130_fd_sc_hd__xor2_1
XTAP_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$576 U$$711/B1 U$$578/A2 U$$578/A1 U$$578/B2 VGND VGND VPWR VPWR U$$577/A sky130_fd_sc_hd__a22o_1
XFILLER_44_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$587 U$$587/A U$$607/B VGND VGND VPWR VPWR U$$587/X sky130_fd_sc_hd__xor2_1
XFILLER_204_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$598 U$$598/A1 U$$616/A2 U$$598/B1 U$$616/B2 VGND VGND VPWR VPWR U$$599/A sky130_fd_sc_hd__a22o_1
XFILLER_60_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_528 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1410 input25/X VGND VGND VPWR VPWR U$$2178/B sky130_fd_sc_hd__buf_6
Xrepeater1421 U$$1912/B VGND VGND VPWR VPWR U$$1870/B sky130_fd_sc_hd__buf_6
XFILLER_67_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1432 U$$1751/B VGND VGND VPWR VPWR U$$1679/B sky130_fd_sc_hd__buf_8
XFILLER_126_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1443 U$$1608/B VGND VGND VPWR VPWR U$$1592/B sky130_fd_sc_hd__buf_8
XFILLER_153_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1454 U$$1507/A VGND VGND VPWR VPWR U$$1499/B sky130_fd_sc_hd__buf_6
XFILLER_67_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_88_5 dadda_fa_2_88_5/A dadda_fa_2_88_5/B dadda_fa_2_88_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_89_2/A dadda_fa_4_88_0/A sky130_fd_sc_hd__fa_2
Xrepeater1465 U$$983/A1 VGND VGND VPWR VPWR U$$1666/B1 sky130_fd_sc_hd__buf_4
Xrepeater1476 U$$4269/A1 VGND VGND VPWR VPWR U$$3447/A1 sky130_fd_sc_hd__buf_6
XFILLER_193_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1487 U$$431/A1 VGND VGND VPWR VPWR U$$4404/A1 sky130_fd_sc_hd__buf_12
XFILLER_119_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1498 U$$954/A1 VGND VGND VPWR VPWR U$$678/B1 sky130_fd_sc_hd__buf_4
XFILLER_99_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_31_1 U$$468/X U$$601/X U$$734/X VGND VGND VPWR VPWR dadda_fa_3_32_1/A
+ dadda_fa_3_31_3/A sky130_fd_sc_hd__fa_1
XFILLER_36_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_24_0 U$$55/X U$$188/X U$$321/X VGND VGND VPWR VPWR dadda_fa_3_25_3/A dadda_fa_3_24_3/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_211_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1260 U$$1260/A U$$1330/B VGND VGND VPWR VPWR U$$1260/X sky130_fd_sc_hd__xor2_1
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1271 U$$721/B1 U$$1271/A2 U$$999/A1 U$$1271/B2 VGND VGND VPWR VPWR U$$1272/A sky130_fd_sc_hd__a22o_1
XU$$1282 U$$1282/A U$$1286/B VGND VGND VPWR VPWR U$$1282/X sky130_fd_sc_hd__xor2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1293 U$$60/A1 U$$1337/A2 U$$62/A1 U$$1337/B2 VGND VGND VPWR VPWR U$$1294/A sky130_fd_sc_hd__a22o_1
XFILLER_202_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_118_1 dadda_fa_5_118_1/A dadda_fa_5_118_1/B dadda_ha_4_118_2/SUM VGND
+ VGND VPWR VPWR dadda_fa_6_119_0/B dadda_fa_7_118_0/A sky130_fd_sc_hd__fa_1
Xdadda_ha_1_84_6 U$$3766/X U$$3899/X VGND VGND VPWR VPWR dadda_fa_2_85_4/A dadda_fa_3_84_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_83_4 U$$2966/X U$$3099/X U$$3232/X VGND VGND VPWR VPWR dadda_fa_2_84_3/A
+ dadda_fa_2_83_5/B sky130_fd_sc_hd__fa_1
XFILLER_172_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_76_3 U$$2686/X U$$2819/X U$$2952/X VGND VGND VPWR VPWR dadda_fa_2_77_1/B
+ dadda_fa_2_76_4/B sky130_fd_sc_hd__fa_1
XFILLER_113_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_53_2 dadda_fa_4_53_2/A dadda_fa_4_53_2/B dadda_fa_4_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_54_0/CIN dadda_fa_5_53_1/CIN sky130_fd_sc_hd__fa_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_2 U$$3204/X U$$3337/X U$$3470/X VGND VGND VPWR VPWR dadda_fa_2_70_1/A
+ dadda_fa_2_69_4/A sky130_fd_sc_hd__fa_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_46_1 dadda_fa_4_46_1/A dadda_fa_4_46_1/B dadda_fa_4_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/B dadda_fa_5_46_1/B sky130_fd_sc_hd__fa_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_23_0 dadda_fa_7_23_0/A dadda_fa_7_23_0/B dadda_fa_7_23_0/CIN VGND VGND
+ VPWR VPWR _320_/D _191_/D sky130_fd_sc_hd__fa_2
XFILLER_22_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_39_0 dadda_fa_4_39_0/A dadda_fa_4_39_0/B dadda_fa_4_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/A dadda_fa_5_39_1/A sky130_fd_sc_hd__fa_1
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _199_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_216 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_227 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_249 U$$3293/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ _360_/CLK _360_/D VGND VGND VPWR VPWR _360_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_291_ _420_/CLK _291_/D VGND VGND VPWR VPWR _291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_336 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_71_2 U$$1346/X U$$1479/X U$$1612/X VGND VGND VPWR VPWR dadda_fa_1_72_7/B
+ dadda_fa_1_71_8/CIN sky130_fd_sc_hd__fa_1
XTAP_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_64_1 U$$534/X U$$667/X U$$800/X VGND VGND VPWR VPWR dadda_fa_1_65_5/CIN
+ dadda_fa_1_64_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_41_0 dadda_fa_3_41_0/A dadda_fa_3_41_0/B dadda_fa_3_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_0/B dadda_fa_4_41_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1028 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_57_0 U$$121/X U$$254/X U$$387/X VGND VGND VPWR VPWR dadda_fa_1_58_7/A
+ dadda_fa_1_57_8/B sky130_fd_sc_hd__fa_1
XTAP_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$490 final_adder.U$$494/B final_adder.U$$490/B VGND VGND VPWR VPWR
+ final_adder.U$$614/B sky130_fd_sc_hd__and2_1
XTAP_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$340 U$$66/A1 U$$340/A2 U$$68/A1 U$$340/B2 VGND VGND VPWR VPWR U$$341/A sky130_fd_sc_hd__a22o_1
XTAP_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$351 U$$351/A U$$351/B VGND VGND VPWR VPWR U$$351/X sky130_fd_sc_hd__xor2_1
XTAP_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$362 U$$88/A1 U$$396/A2 U$$90/A1 U$$396/B2 VGND VGND VPWR VPWR U$$363/A sky130_fd_sc_hd__a22o_1
XFILLER_32_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$373 U$$373/A U$$377/B VGND VGND VPWR VPWR U$$373/X sky130_fd_sc_hd__xor2_1
XFILLER_205_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$384 U$$384/A1 U$$394/A2 U$$384/B1 U$$394/B2 VGND VGND VPWR VPWR U$$385/A sky130_fd_sc_hd__a22o_1
XU$$395 U$$395/A U$$395/B VGND VGND VPWR VPWR U$$395/X sky130_fd_sc_hd__xor2_1
XFILLER_60_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_93_3 U$$4050/X U$$4183/X U$$4316/X VGND VGND VPWR VPWR dadda_fa_3_94_1/B
+ dadda_fa_3_93_3/B sky130_fd_sc_hd__fa_1
XFILLER_114_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1240 input58/X VGND VGND VPWR VPWR U$$4243/B sky130_fd_sc_hd__buf_4
Xrepeater1251 U$$4100/B VGND VGND VPWR VPWR U$$4080/B sky130_fd_sc_hd__buf_6
XFILLER_160_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_86_2 input241/X dadda_fa_2_86_2/B dadda_fa_2_86_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_87_1/A dadda_fa_3_86_3/A sky130_fd_sc_hd__fa_1
XFILLER_5_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1262 U$$3875/B VGND VGND VPWR VPWR U$$3879/B sky130_fd_sc_hd__buf_6
XFILLER_99_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1273 U$$3834/B VGND VGND VPWR VPWR U$$3826/B sky130_fd_sc_hd__buf_8
XFILLER_113_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1284 input5/X VGND VGND VPWR VPWR U$$959/A sky130_fd_sc_hd__buf_4
XFILLER_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1295 U$$3490/B VGND VGND VPWR VPWR U$$3528/B sky130_fd_sc_hd__buf_8
Xdadda_fa_5_63_1 dadda_fa_5_63_1/A dadda_fa_5_63_1/B dadda_fa_5_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_64_0/B dadda_fa_7_63_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_79_1 dadda_fa_2_79_1/A dadda_fa_2_79_1/B dadda_fa_2_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_0/CIN dadda_fa_3_79_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_778 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_56_0 dadda_fa_5_56_0/A dadda_fa_5_56_0/B dadda_fa_5_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_57_0/A dadda_fa_6_56_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1367_1715 VGND VGND VPWR VPWR U$$1367_1715/HI U$$1367/B1 sky130_fd_sc_hd__conb_1
XFILLER_171_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1038 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_55_8 dadda_fa_1_55_8/A dadda_fa_1_55_8/B dadda_fa_1_55_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_56_3/A dadda_fa_3_55_0/A sky130_fd_sc_hd__fa_1
XFILLER_28_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_102_0 dadda_fa_2_102_0/A U$$2738/X U$$2871/X VGND VGND VPWR VPWR dadda_fa_3_103_2/A
+ dadda_fa_3_102_3/A sky130_fd_sc_hd__fa_1
XFILLER_63_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1090 U$$1090/A U$$1095/A VGND VGND VPWR VPWR U$$1090/X sky130_fd_sc_hd__xor2_1
XFILLER_10_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2326_1730 VGND VGND VPWR VPWR U$$2326_1730/HI U$$2326/B1 sky130_fd_sc_hd__conb_1
XFILLER_191_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_81_1 U$$1632/X U$$1765/X U$$1898/X VGND VGND VPWR VPWR dadda_fa_2_82_1/B
+ dadda_fa_2_81_4/A sky130_fd_sc_hd__fa_1
XFILLER_176_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_74_0 U$$1751/X U$$1884/X U$$2017/X VGND VGND VPWR VPWR dadda_fa_2_75_0/B
+ dadda_fa_2_74_3/B sky130_fd_sc_hd__fa_1
XFILLER_137_1088 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3409 U$$3409/A U$$3424/A VGND VGND VPWR VPWR U$$3409/X sky130_fd_sc_hd__xor2_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2708 U$$2708/A U$$2710/B VGND VGND VPWR VPWR U$$2708/X sky130_fd_sc_hd__xor2_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2719 U$$4361/B1 U$$2737/A2 U$$4228/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2720/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_412_ _412_/CLK _412_/D VGND VGND VPWR VPWR _412_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_502 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_343_ _351_/CLK _343_/D VGND VGND VPWR VPWR _343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_274_ _407_/CLK _274_/D VGND VGND VPWR VPWR _274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_96_1 dadda_fa_3_96_1/A dadda_fa_3_96_1/B dadda_fa_3_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_0/CIN dadda_fa_4_96_2/A sky130_fd_sc_hd__fa_1
XFILLER_143_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_73_0 dadda_fa_6_73_0/A dadda_fa_6_73_0/B dadda_fa_6_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_74_0/B dadda_fa_7_73_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_136_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_89_0 dadda_fa_3_89_0/A dadda_fa_3_89_0/B dadda_fa_3_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_0/B dadda_fa_4_89_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_190_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater907 U$$3648/B1 VGND VGND VPWR VPWR U$$2691/A1 sky130_fd_sc_hd__buf_6
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater918 input98/X VGND VGND VPWR VPWR U$$3713/A1 sky130_fd_sc_hd__buf_4
XFILLER_204_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater929 U$$4055/B1 VGND VGND VPWR VPWR U$$2550/A1 sky130_fd_sc_hd__buf_6
XFILLER_77_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3910 input91/X U$$3970/A2 input92/X U$$3970/B2 VGND VGND VPWR VPWR U$$3911/A sky130_fd_sc_hd__a22o_1
XFILLER_209_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3921 U$$3921/A U$$3927/B VGND VGND VPWR VPWR U$$3921/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_118_0 dadda_fa_4_118_0/A U$$3834/X U$$3967/X VGND VGND VPWR VPWR dadda_fa_5_119_0/B
+ dadda_fa_5_118_1/A sky130_fd_sc_hd__fa_1
XFILLER_94_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3932 U$$4343/A1 U$$3946/A2 U$$4343/B1 U$$3946/B2 VGND VGND VPWR VPWR U$$3933/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3943 U$$3943/A U$$3947/B VGND VGND VPWR VPWR U$$3943/X sky130_fd_sc_hd__xor2_1
XTAP_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3954 input115/X U$$3968/A2 U$$4504/A1 U$$3968/B2 VGND VGND VPWR VPWR U$$3955/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_5_5_0 U$$17/X U$$150/X VGND VGND VPWR VPWR dadda_fa_6_6_0/B dadda_fa_7_5_0/A
+ sky130_fd_sc_hd__ha_1
XU$$3965 U$$3965/A U$$3972/A VGND VGND VPWR VPWR U$$3965/X sky130_fd_sc_hd__xor2_1
XFILLER_24_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3976 U$$4109/A U$$3976/B VGND VGND VPWR VPWR U$$3976/X sky130_fd_sc_hd__and2_1
XTAP_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3987 U$$4398/A1 U$$4011/A2 U$$3987/B1 U$$4011/B2 VGND VGND VPWR VPWR U$$3988/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3998 U$$3998/A U$$4036/B VGND VGND VPWR VPWR U$$3998/X sky130_fd_sc_hd__xor2_1
XFILLER_80_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$170 U$$170/A U$$176/B VGND VGND VPWR VPWR U$$170/X sky130_fd_sc_hd__xor2_1
XFILLER_73_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$181 U$$44/A1 U$$209/A2 U$$46/A1 U$$209/B2 VGND VGND VPWR VPWR U$$182/A sky130_fd_sc_hd__a22o_1
XU$$192 U$$192/A U$$218/B VGND VGND VPWR VPWR U$$192/X sky130_fd_sc_hd__xor2_1
XFILLER_205_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_91_0 U$$3115/X U$$3248/X U$$3381/X VGND VGND VPWR VPWR dadda_fa_3_92_0/B
+ dadda_fa_3_91_2/B sky130_fd_sc_hd__fa_1
XFILLER_145_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1070 U$$4162/B1 VGND VGND VPWR VPWR U$$4438/A1 sky130_fd_sc_hd__buf_6
Xoutput267 output267/A VGND VGND VPWR VPWR o[109] sky130_fd_sc_hd__buf_2
XFILLER_173_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1081 input79/X VGND VGND VPWR VPWR U$$4162/A1 sky130_fd_sc_hd__buf_6
Xrepeater1092 U$$4293/B1 VGND VGND VPWR VPWR U$$4432/A1 sky130_fd_sc_hd__buf_4
XFILLER_114_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput278 output278/A VGND VGND VPWR VPWR o[119] sky130_fd_sc_hd__buf_2
XFILLER_102_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput289 output289/A VGND VGND VPWR VPWR o[13] sky130_fd_sc_hd__buf_2
XFILLER_47_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_1_47_6 U$$2495/X U$$2628/X VGND VGND VPWR VPWR dadda_fa_2_48_3/B dadda_fa_3_47_0/A
+ sky130_fd_sc_hd__ha_1
XU$$1230_1712 VGND VGND VPWR VPWR U$$1230_1712/HI U$$1230/B1 sky130_fd_sc_hd__conb_1
XFILLER_101_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_60_6 input213/X dadda_fa_1_60_6/B dadda_fa_1_60_6/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_61_2/B dadda_fa_2_60_5/B sky130_fd_sc_hd__fa_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_5 U$$2374/X U$$2507/X U$$2640/X VGND VGND VPWR VPWR dadda_fa_2_54_2/A
+ dadda_fa_2_53_5/A sky130_fd_sc_hd__fa_1
XFILLER_210_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_46_4 U$$1695/X U$$1828/X U$$1961/X VGND VGND VPWR VPWR dadda_fa_2_47_3/A
+ dadda_fa_2_46_5/B sky130_fd_sc_hd__fa_1
XFILLER_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_16_2 dadda_fa_4_16_2/A dadda_fa_4_16_2/B dadda_ha_3_16_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_17_0/CIN dadda_fa_5_16_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_24_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_90_0 dadda_fa_7_90_0/A dadda_fa_7_90_0/B dadda_fa_7_90_0/CIN VGND VGND
+ VPWR VPWR _387_/D _258_/D sky130_fd_sc_hd__fa_1
XFILLER_183_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1108 final_adder.U$$170/A final_adder.U$$879/X VGND VGND VPWR VPWR
+ output367/A sky130_fd_sc_hd__xor2_1
XFILLER_177_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$1119 final_adder.U$$160/B final_adder.U$$931/X VGND VGND VPWR VPWR
+ output379/A sky130_fd_sc_hd__xor2_1
XFILLER_20_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3206 U$$3206/A U$$3244/B VGND VGND VPWR VPWR U$$3206/X sky130_fd_sc_hd__xor2_1
XFILLER_74_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3217 U$$4450/A1 U$$3255/A2 U$$4452/A1 U$$3255/B2 VGND VGND VPWR VPWR U$$3218/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3228 U$$3228/A U$$3228/B VGND VGND VPWR VPWR U$$3228/X sky130_fd_sc_hd__xor2_1
XFILLER_189_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3239 U$$3376/A1 U$$3241/A2 U$$3378/A1 U$$3241/B2 VGND VGND VPWR VPWR U$$3240/A
+ sky130_fd_sc_hd__a22o_1
XU$$2505 U$$2505/A U$$2597/B VGND VGND VPWR VPWR U$$2505/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2516 U$$50/A1 U$$2542/A2 U$$3612/B1 U$$2542/B2 VGND VGND VPWR VPWR U$$2517/A sky130_fd_sc_hd__a22o_1
XFILLER_185_1137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2527 U$$2527/A U$$2577/B VGND VGND VPWR VPWR U$$2527/X sky130_fd_sc_hd__xor2_1
XFILLER_64_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2538 U$$2810/B1 U$$2558/A2 U$$3499/A1 U$$2558/B2 VGND VGND VPWR VPWR U$$2539/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1804 U$$1804/A U$$1840/B VGND VGND VPWR VPWR U$$1804/X sky130_fd_sc_hd__xor2_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2549 U$$2549/A U$$2601/B VGND VGND VPWR VPWR U$$2549/X sky130_fd_sc_hd__xor2_1
XU$$1815 U$$993/A1 U$$1819/A2 U$$993/B1 U$$1819/B2 VGND VGND VPWR VPWR U$$1816/A sky130_fd_sc_hd__a22o_1
XFILLER_61_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1826 U$$1826/A U$$1878/B VGND VGND VPWR VPWR U$$1826/X sky130_fd_sc_hd__xor2_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1837 U$$3481/A1 U$$1839/A2 U$$3618/B1 U$$1839/B2 VGND VGND VPWR VPWR U$$1838/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1848 U$$1848/A U$$1880/B VGND VGND VPWR VPWR U$$1848/X sky130_fd_sc_hd__xor2_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1859 U$$763/A1 U$$1869/A2 U$$763/B1 U$$1869/B2 VGND VGND VPWR VPWR U$$1860/A sky130_fd_sc_hd__a22o_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_326_ _326_/CLK _326_/D VGND VGND VPWR VPWR _326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_257_ _387_/CLK _257_/D VGND VGND VPWR VPWR _257_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_188_ _329_/CLK _188_/D VGND VGND VPWR VPWR _188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_70_5 dadda_fa_2_70_5/A dadda_fa_2_70_5/B dadda_fa_2_70_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_2/A dadda_fa_4_70_0/A sky130_fd_sc_hd__fa_1
XU$$4390_1771 VGND VGND VPWR VPWR U$$4390_1771/HI U$$4390/A1 sky130_fd_sc_hd__conb_1
XFILLER_42_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_63_4 dadda_fa_2_63_4/A dadda_fa_2_63_4/B dadda_fa_2_63_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_1/CIN dadda_fa_3_63_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater704 U$$3970/B2 VGND VGND VPWR VPWR U$$3874/B2 sky130_fd_sc_hd__clkbuf_8
Xrepeater715 U$$3773/B2 VGND VGND VPWR VPWR U$$3739/B2 sky130_fd_sc_hd__buf_4
XFILLER_78_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater726 U$$3430/X VGND VGND VPWR VPWR U$$3503/B2 sky130_fd_sc_hd__buf_4
Xrepeater737 U$$3416/B2 VGND VGND VPWR VPWR U$$3422/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_56_3 dadda_fa_2_56_3/A dadda_fa_2_56_3/B dadda_fa_2_56_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/B dadda_fa_3_56_3/B sky130_fd_sc_hd__fa_1
XFILLER_42_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater748 U$$3255/B2 VGND VGND VPWR VPWR U$$3285/B2 sky130_fd_sc_hd__buf_6
XU$$4430 U$$4430/A1 U$$4388/X U$$4432/A1 U$$4430/B2 VGND VGND VPWR VPWR U$$4431/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater759 U$$2985/B2 VGND VGND VPWR VPWR U$$3011/B2 sky130_fd_sc_hd__buf_6
XU$$4441 U$$4441/A U$$4441/B VGND VGND VPWR VPWR U$$4441/X sky130_fd_sc_hd__xor2_1
XU$$4452 U$$4452/A1 U$$4388/X U$$4454/A1 U$$4476/B2 VGND VGND VPWR VPWR U$$4453/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_49_2 dadda_fa_2_49_2/A dadda_fa_2_49_2/B dadda_fa_2_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/A dadda_fa_3_49_3/A sky130_fd_sc_hd__fa_1
XU$$4463 U$$4463/A U$$4463/B VGND VGND VPWR VPWR U$$4463/X sky130_fd_sc_hd__xor2_1
XFILLER_42_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4474 input100/X U$$4388/X input101/X U$$4486/B2 VGND VGND VPWR VPWR U$$4475/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4485 U$$4485/A U$$4485/B VGND VGND VPWR VPWR U$$4485/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_26_1 dadda_fa_5_26_1/A dadda_fa_5_26_1/B dadda_fa_5_26_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_27_0/B dadda_fa_7_26_0/A sky130_fd_sc_hd__fa_2
XU$$3740 U$$3740/A U$$3740/B VGND VGND VPWR VPWR U$$3740/X sky130_fd_sc_hd__xor2_1
XU$$4496 U$$4496/A1 U$$4388/X U$$4498/A1 U$$4498/B2 VGND VGND VPWR VPWR U$$4497/A
+ sky130_fd_sc_hd__a22o_1
XU$$3751 input79/X U$$3793/A2 input80/X U$$3793/B2 VGND VGND VPWR VPWR U$$3752/A sky130_fd_sc_hd__a22o_1
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3762 U$$3762/A U$$3836/A VGND VGND VPWR VPWR U$$3762/X sky130_fd_sc_hd__xor2_1
XFILLER_25_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3773 U$$3908/B1 U$$3773/A2 U$$3775/A1 U$$3773/B2 VGND VGND VPWR VPWR U$$3774/A
+ sky130_fd_sc_hd__a22o_1
XU$$3784 U$$3784/A U$$3814/B VGND VGND VPWR VPWR U$$3784/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_19_0 dadda_fa_5_19_0/A dadda_fa_5_19_0/B dadda_fa_5_19_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_20_0/A dadda_fa_6_19_0/CIN sky130_fd_sc_hd__fa_1
XU$$3795 U$$4343/A1 U$$3813/A2 U$$4343/B1 U$$3813/B2 VGND VGND VPWR VPWR U$$3796/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_280 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_100_1 dadda_fa_5_100_1/A dadda_fa_5_100_1/B dadda_fa_5_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_101_0/B dadda_fa_7_100_0/A sky130_fd_sc_hd__fa_1
XU$$4473_1813 VGND VGND VPWR VPWR U$$4473_1813/HI U$$4473/B sky130_fd_sc_hd__conb_1
XFILLER_106_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_4_122_0 dadda_ha_4_122_0/A U$$4108/X VGND VGND VPWR VPWR dadda_fa_5_123_1/CIN
+ dadda_ha_4_122_0/SUM sky130_fd_sc_hd__ha_1
XFILLER_133_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_38_2 U$$881/X U$$1014/X VGND VGND VPWR VPWR dadda_fa_2_39_5/A dadda_fa_3_38_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_102_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_51_2 U$$907/X U$$1040/X U$$1173/X VGND VGND VPWR VPWR dadda_fa_2_52_1/A
+ dadda_fa_2_51_4/A sky130_fd_sc_hd__fa_1
XU$$906 U$$84/A1 U$$906/A2 U$$84/B1 U$$906/B2 VGND VGND VPWR VPWR U$$907/A sky130_fd_sc_hd__a22o_1
XU$$917 U$$917/A U$$958/A VGND VGND VPWR VPWR U$$917/X sky130_fd_sc_hd__xor2_1
XFILLER_56_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$928 U$$928/A1 U$$938/A2 U$$930/A1 U$$938/B2 VGND VGND VPWR VPWR U$$929/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_44_1 U$$494/X U$$627/X U$$760/X VGND VGND VPWR VPWR dadda_fa_2_45_2/CIN
+ dadda_fa_2_44_4/CIN sky130_fd_sc_hd__fa_1
XU$$939 U$$939/A U$$959/A VGND VGND VPWR VPWR U$$939/X sky130_fd_sc_hd__xor2_1
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_21_0 input170/X dadda_fa_4_21_0/B dadda_fa_4_21_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_5_22_0/A dadda_fa_5_21_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_37_0 U$$81/X U$$214/X U$$347/X VGND VGND VPWR VPWR dadda_fa_2_38_4/CIN
+ dadda_fa_2_37_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_5_126_0_1876 VGND VGND VPWR VPWR dadda_ha_5_126_0/A dadda_ha_5_126_0_1876/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_180_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_73_3 dadda_fa_3_73_3/A dadda_fa_3_73_3/B dadda_fa_3_73_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_74_1/B dadda_fa_4_73_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_1106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_66_2 dadda_fa_3_66_2/A dadda_fa_3_66_2/B dadda_fa_3_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_1/A dadda_fa_4_66_2/B sky130_fd_sc_hd__fa_1
XFILLER_152_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_59_1 dadda_fa_3_59_1/A dadda_fa_3_59_1/B dadda_fa_3_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_0/CIN dadda_fa_4_59_2/A sky130_fd_sc_hd__fa_1
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_36_0 dadda_fa_6_36_0/A dadda_fa_6_36_0/B dadda_fa_6_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_37_0/B dadda_fa_7_36_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_8_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3003 U$$3551/A1 U$$3011/A2 input121/X U$$3011/B2 VGND VGND VPWR VPWR U$$3004/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3014 input38/X VGND VGND VPWR VPWR U$$3014/Y sky130_fd_sc_hd__inv_1
XFILLER_93_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3025 U$$3025/A U$$3075/B VGND VGND VPWR VPWR U$$3025/X sky130_fd_sc_hd__xor2_1
XU$$3036 U$$842/B1 U$$3124/A2 U$$24/A1 U$$3124/B2 VGND VGND VPWR VPWR U$$3037/A sky130_fd_sc_hd__a22o_1
XU$$2302 U$$2711/B1 U$$2302/A2 U$$934/A1 U$$2302/B2 VGND VGND VPWR VPWR U$$2303/A
+ sky130_fd_sc_hd__a22o_1
XU$$3047 U$$3047/A U$$3125/B VGND VGND VPWR VPWR U$$3047/X sky130_fd_sc_hd__xor2_1
XU$$3058 U$$3058/A1 U$$3060/A2 U$$3606/B1 U$$3060/B2 VGND VGND VPWR VPWR U$$3059/A
+ sky130_fd_sc_hd__a22o_1
XU$$2313 U$$2313/A input27/X VGND VGND VPWR VPWR U$$2313/X sky130_fd_sc_hd__xor2_1
XFILLER_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2324 U$$2324/A1 U$$2326/A2 U$$956/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2325/A
+ sky130_fd_sc_hd__a22o_1
XU$$3069 U$$3069/A U$$3077/B VGND VGND VPWR VPWR U$$3069/X sky130_fd_sc_hd__xor2_1
XFILLER_90_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2335 U$$2335/A1 U$$2417/A2 U$$2609/B1 U$$2417/B2 VGND VGND VPWR VPWR U$$2336/A
+ sky130_fd_sc_hd__a22o_1
XU$$1601 U$$3108/A1 U$$1607/A2 U$$3108/B1 U$$1607/B2 VGND VGND VPWR VPWR U$$1602/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2346 U$$2346/A U$$2360/B VGND VGND VPWR VPWR U$$2346/X sky130_fd_sc_hd__xor2_1
XFILLER_201_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2357 U$$3453/A1 U$$2403/A2 U$$2357/B1 U$$2403/B2 VGND VGND VPWR VPWR U$$2358/A
+ sky130_fd_sc_hd__a22o_1
XU$$1612 U$$1612/A U$$1628/B VGND VGND VPWR VPWR U$$1612/X sky130_fd_sc_hd__xor2_1
XU$$1623 U$$527/A1 U$$1635/A2 U$$527/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1624/A sky130_fd_sc_hd__a22o_1
XU$$2368 U$$2368/A U$$2380/B VGND VGND VPWR VPWR U$$2368/X sky130_fd_sc_hd__xor2_1
XU$$2379 U$$3749/A1 U$$2463/A2 U$$3749/B1 U$$2463/B2 VGND VGND VPWR VPWR U$$2380/A
+ sky130_fd_sc_hd__a22o_1
XU$$1634 U$$1634/A U$$1638/B VGND VGND VPWR VPWR U$$1634/X sky130_fd_sc_hd__xor2_1
XFILLER_90_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1645 input17/X VGND VGND VPWR VPWR U$$1647/B sky130_fd_sc_hd__inv_1
XFILLER_76_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1656 U$$2065/B1 U$$1688/A2 U$$2343/A1 U$$1688/B2 VGND VGND VPWR VPWR U$$1657/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1667 U$$1667/A U$$1679/B VGND VGND VPWR VPWR U$$1667/X sky130_fd_sc_hd__xor2_1
XFILLER_199_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1678 U$$993/A1 U$$1696/A2 U$$993/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1679/A sky130_fd_sc_hd__a22o_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1689 U$$1689/A U$$1689/B VGND VGND VPWR VPWR U$$1689/X sky130_fd_sc_hd__xor2_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_309_ _314_/CLK _309_/D VGND VGND VPWR VPWR _309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_109_0 dadda_fa_7_109_0/A dadda_fa_7_109_0/B dadda_fa_7_109_0/CIN VGND
+ VGND VPWR VPWR _406_/D _277_/D sky130_fd_sc_hd__fa_1
XFILLER_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_61_1 dadda_fa_2_61_1/A dadda_fa_2_61_1/B dadda_fa_2_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_0/CIN dadda_fa_3_61_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater501 U$$3155/X VGND VGND VPWR VPWR U$$3241/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$308 final_adder.U$$310/B final_adder.U$$308/B VGND VGND VPWR VPWR
+ final_adder.U$$434/B sky130_fd_sc_hd__and2_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater512 U$$2985/A2 VGND VGND VPWR VPWR U$$3011/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$319 final_adder.U$$318/B final_adder.U$$193/X final_adder.U$$191/X
+ VGND VGND VPWR VPWR final_adder.U$$319/X sky130_fd_sc_hd__a21o_1
Xrepeater523 U$$366/A2 VGND VGND VPWR VPWR U$$378/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_54_0 dadda_fa_2_54_0/A dadda_fa_2_54_0/B dadda_fa_2_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_0/B dadda_fa_3_54_2/B sky130_fd_sc_hd__fa_1
XFILLER_38_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater534 U$$2844/A2 VGND VGND VPWR VPWR U$$2828/A2 sky130_fd_sc_hd__buf_6
Xrepeater545 U$$2588/A2 VGND VGND VPWR VPWR U$$2600/A2 sky130_fd_sc_hd__buf_4
Xrepeater556 U$$2459/A2 VGND VGND VPWR VPWR U$$2463/A2 sky130_fd_sc_hd__buf_4
Xrepeater567 U$$2091/A2 VGND VGND VPWR VPWR U$$2093/A2 sky130_fd_sc_hd__buf_4
XU$$4260 U$$4260/A U$$4278/B VGND VGND VPWR VPWR U$$4260/X sky130_fd_sc_hd__xor2_1
XFILLER_66_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater578 U$$2022/A2 VGND VGND VPWR VPWR U$$2016/A2 sky130_fd_sc_hd__buf_6
Xrepeater589 U$$1913/A2 VGND VGND VPWR VPWR U$$1877/A2 sky130_fd_sc_hd__buf_8
XU$$4271 U$$4408/A1 U$$4275/A2 U$$4408/B1 U$$4275/B2 VGND VGND VPWR VPWR U$$4272/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3559_1750 VGND VGND VPWR VPWR U$$3559_1750/HI U$$3559/B1 sky130_fd_sc_hd__conb_1
XU$$4282 U$$4282/A U$$4330/B VGND VGND VPWR VPWR U$$4282/X sky130_fd_sc_hd__xor2_1
XU$$4293 input75/X U$$4297/A2 U$$4293/B1 U$$4297/B2 VGND VGND VPWR VPWR U$$4294/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3570 U$$3979/B1 U$$3612/A2 U$$832/A1 U$$3612/B2 VGND VGND VPWR VPWR U$$3571/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3581 U$$3581/A U$$3609/B VGND VGND VPWR VPWR U$$3581/X sky130_fd_sc_hd__xor2_1
XU$$3592 U$$3727/B1 U$$3606/A2 U$$4005/A1 U$$3606/B2 VGND VGND VPWR VPWR U$$3593/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_991 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_8_0 U$$289/X U$$422/X U$$555/X VGND VGND VPWR VPWR dadda_fa_6_9_0/A dadda_fa_6_8_0/CIN
+ sky130_fd_sc_hd__fa_1
XU$$2880 input38/X U$$2880/B VGND VGND VPWR VPWR U$$2880/X sky130_fd_sc_hd__and2_1
XU$$2891 U$$4398/A1 U$$2921/A2 U$$3987/B1 U$$2921/B2 VGND VGND VPWR VPWR U$$2892/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_83_2 dadda_fa_4_83_2/A dadda_fa_4_83_2/B dadda_fa_4_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_84_0/CIN dadda_fa_5_83_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_76_1 dadda_fa_4_76_1/A dadda_fa_4_76_1/B dadda_fa_4_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/B dadda_fa_5_76_1/B sky130_fd_sc_hd__fa_1
XFILLER_161_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_53_0 dadda_fa_7_53_0/A dadda_fa_7_53_0/B dadda_fa_7_53_0/CIN VGND VGND
+ VPWR VPWR _350_/D _221_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_69_0 dadda_fa_4_69_0/A dadda_fa_4_69_0/B dadda_fa_4_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/A dadda_fa_5_69_1/A sky130_fd_sc_hd__fa_1
XFILLER_88_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$831 final_adder.U$$798/A final_adder.U$$381/X final_adder.U$$719/X
+ VGND VGND VPWR VPWR final_adder.U$$831/X sky130_fd_sc_hd__a21o_1
XTAP_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$853 final_adder.U$$756/X final_adder.U$$821/X final_adder.U$$757/X
+ VGND VGND VPWR VPWR final_adder.U$$853/X sky130_fd_sc_hd__a21o_2
XFILLER_25_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$703 U$$703/A1 U$$711/A2 U$$979/A1 U$$711/B2 VGND VGND VPWR VPWR U$$704/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$875 final_adder.U$$778/X final_adder.U$$731/X final_adder.U$$779/X
+ VGND VGND VPWR VPWR final_adder.U$$875/X sky130_fd_sc_hd__a21o_1
XU$$714 U$$714/A U$$740/B VGND VGND VPWR VPWR U$$714/X sky130_fd_sc_hd__xor2_1
XFILLER_99_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$725 U$$860/B1 U$$759/A2 U$$727/A1 U$$759/B2 VGND VGND VPWR VPWR U$$726/A sky130_fd_sc_hd__a22o_1
XFILLER_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$897 final_adder.U$$800/X final_adder.U$$255/X final_adder.U$$801/X
+ VGND VGND VPWR VPWR final_adder.U$$897/X sky130_fd_sc_hd__a21o_1
XU$$736 U$$736/A U$$770/B VGND VGND VPWR VPWR U$$736/X sky130_fd_sc_hd__xor2_1
XU$$747 U$$882/B1 U$$749/A2 U$$64/A1 U$$749/B2 VGND VGND VPWR VPWR U$$748/A sky130_fd_sc_hd__a22o_1
XFILLER_83_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$758 U$$758/A U$$796/B VGND VGND VPWR VPWR U$$758/X sky130_fd_sc_hd__xor2_1
XFILLER_44_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$769 U$$84/A1 U$$793/A2 U$$84/B1 U$$793/B2 VGND VGND VPWR VPWR U$$770/A sky130_fd_sc_hd__a22o_1
XFILLER_72_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1603 U$$3944/B1 VGND VGND VPWR VPWR U$$521/A1 sky130_fd_sc_hd__buf_4
XFILLER_32_1187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_8 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1614 U$$2848/A1 VGND VGND VPWR VPWR U$$930/A1 sky130_fd_sc_hd__buf_12
Xrepeater1625 U$$1366/B VGND VGND VPWR VPWR U$$1316/B sky130_fd_sc_hd__buf_6
XFILLER_4_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1636 input109/X VGND VGND VPWR VPWR U$$3852/A1 sky130_fd_sc_hd__buf_4
Xrepeater1647 U$$4488/A1 VGND VGND VPWR VPWR U$$3801/B1 sky130_fd_sc_hd__buf_4
XFILLER_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1658 U$$3116/A1 VGND VGND VPWR VPWR U$$2292/B1 sky130_fd_sc_hd__buf_6
XFILLER_125_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1669 input104/X VGND VGND VPWR VPWR U$$4343/B1 sky130_fd_sc_hd__buf_4
XFILLER_180_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_71_0 dadda_fa_3_71_0/A dadda_fa_3_71_0/B dadda_fa_3_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_0/B dadda_fa_4_71_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1097 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2110 U$$2110/A U$$2114/B VGND VGND VPWR VPWR U$$2110/X sky130_fd_sc_hd__xor2_1
XFILLER_47_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_100_0 dadda_fa_4_100_0/A dadda_fa_4_100_0/B dadda_fa_4_100_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/A dadda_fa_5_100_1/A sky130_fd_sc_hd__fa_1
XFILLER_62_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2121 U$$477/A1 U$$2149/A2 U$$2123/A1 U$$2149/B2 VGND VGND VPWR VPWR U$$2122/A
+ sky130_fd_sc_hd__a22o_1
XU$$2132 U$$2132/A U$$2178/B VGND VGND VPWR VPWR U$$2132/X sky130_fd_sc_hd__xor2_1
XFILLER_35_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2143 U$$2415/B1 U$$2149/A2 U$$2282/A1 U$$2149/B2 VGND VGND VPWR VPWR U$$2144/A
+ sky130_fd_sc_hd__a22o_1
XU$$2154 U$$2154/A U$$2191/A VGND VGND VPWR VPWR U$$2154/X sky130_fd_sc_hd__xor2_1
XU$$1420 U$$461/A1 U$$1470/A2 U$$461/B1 U$$1470/B2 VGND VGND VPWR VPWR U$$1421/A sky130_fd_sc_hd__a22o_1
XU$$2165 U$$2165/A1 U$$2059/X U$$2715/A1 U$$2060/X VGND VGND VPWR VPWR U$$2166/A sky130_fd_sc_hd__a22o_1
XU$$2176 U$$2176/A U$$2178/B VGND VGND VPWR VPWR U$$2176/X sky130_fd_sc_hd__xor2_1
XU$$1431 U$$1431/A U$$1459/B VGND VGND VPWR VPWR U$$1431/X sky130_fd_sc_hd__xor2_1
XU$$1442 U$$2949/A1 U$$1448/A2 U$$74/A1 U$$1448/B2 VGND VGND VPWR VPWR U$$1443/A sky130_fd_sc_hd__a22o_1
XU$$2187 U$$4103/B1 U$$2189/A2 U$$3283/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2188/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2198 U$$2198/A1 U$$2226/A2 U$$2198/B1 U$$2226/B2 VGND VGND VPWR VPWR U$$2199/A
+ sky130_fd_sc_hd__a22o_1
XU$$1453 U$$1453/A U$$1501/B VGND VGND VPWR VPWR U$$1453/X sky130_fd_sc_hd__xor2_1
XFILLER_210_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1464 U$$3108/A1 U$$1470/A2 U$$3108/B1 U$$1470/B2 VGND VGND VPWR VPWR U$$1465/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1475 U$$1475/A U$$1507/A VGND VGND VPWR VPWR U$$1475/X sky130_fd_sc_hd__xor2_1
XFILLER_176_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1486 U$$527/A1 U$$1504/A2 U$$392/A1 U$$1504/B2 VGND VGND VPWR VPWR U$$1487/A sky130_fd_sc_hd__a22o_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1497 U$$1497/A U$$1499/B VGND VGND VPWR VPWR U$$1497/X sky130_fd_sc_hd__xor2_1
XFILLER_124_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2463_1732 VGND VGND VPWR VPWR U$$2463_1732/HI U$$2463/B1 sky130_fd_sc_hd__conb_1
XFILLER_175_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_93_1 dadda_fa_5_93_1/A dadda_fa_5_93_1/B dadda_fa_5_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_94_0/B dadda_fa_7_93_0/A sky130_fd_sc_hd__fa_1
XFILLER_175_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_86_0 dadda_fa_5_86_0/A dadda_fa_5_86_0/B dadda_fa_5_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_87_0/A dadda_fa_6_86_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_190_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_78_7 U$$4020/X U$$4153/X U$$4286/X VGND VGND VPWR VPWR dadda_fa_2_79_2/CIN
+ dadda_fa_2_78_5/CIN sky130_fd_sc_hd__fa_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$105 _401_/Q _273_/Q VGND VGND VPWR VPWR final_adder.U$$151/B1 final_adder.U$$150/B
+ sky130_fd_sc_hd__ha_1
XFILLER_131_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$116 _412_/Q _284_/Q VGND VGND VPWR VPWR final_adder.U$$909/B1 final_adder.U$$138/A
+ sky130_fd_sc_hd__ha_1
XFILLER_85_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$127 _423_/Q _295_/Q VGND VGND VPWR VPWR final_adder.U$$127/COUT final_adder.U$$1151/A
+ sky130_fd_sc_hd__ha_2
XFILLER_170_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$138 final_adder.U$$138/A final_adder.U$$138/B VGND VGND VPWR VPWR
+ final_adder.U$$266/B sky130_fd_sc_hd__and2_1
XFILLER_170_1099 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$149 final_adder.U$$148/B final_adder.U$$919/B1 final_adder.U$$149/B1
+ VGND VGND VPWR VPWR final_adder.U$$149/X sky130_fd_sc_hd__a21o_1
XFILLER_38_451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater386 U$$997/A2 VGND VGND VPWR VPWR U$$999/A2 sky130_fd_sc_hd__buf_4
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater397 U$$950/A2 VGND VGND VPWR VPWR U$$918/A2 sky130_fd_sc_hd__buf_4
XU$$4090 U$$4090/A U$$4110/A VGND VGND VPWR VPWR U$$4090/X sky130_fd_sc_hd__xor2_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_754 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_102_2 dadda_fa_3_102_2/A dadda_fa_3_102_2/B dadda_fa_3_102_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_103_1/A dadda_fa_4_102_2/B sky130_fd_sc_hd__fa_1
XFILLER_134_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput101 b[42] VGND VGND VPWR VPWR input101/X sky130_fd_sc_hd__buf_6
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput112 b[52] VGND VGND VPWR VPWR input112/X sky130_fd_sc_hd__buf_6
XFILLER_103_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput123 b[62] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__buf_6
XFILLER_153_1264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput134 c[104] VGND VGND VPWR VPWR input134/X sky130_fd_sc_hd__buf_4
XFILLER_88_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 c[114] VGND VGND VPWR VPWR input145/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_66_5 U$$2134/X U$$2267/X U$$2400/X VGND VGND VPWR VPWR dadda_fa_1_67_7/A
+ dadda_fa_2_66_0/A sky130_fd_sc_hd__fa_2
Xinput156 c[124] VGND VGND VPWR VPWR input156/X sky130_fd_sc_hd__clkbuf_2
XTAP_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_116_0 dadda_fa_6_116_0/A dadda_fa_6_116_0/B dadda_fa_6_116_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_117_0/B dadda_fa_7_116_0/CIN sky130_fd_sc_hd__fa_1
Xinput167 c[19] VGND VGND VPWR VPWR input167/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput178 c[29] VGND VGND VPWR VPWR input178/X sky130_fd_sc_hd__clkbuf_2
XTAP_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 c[39] VGND VGND VPWR VPWR input189/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$650 final_adder.U$$666/B final_adder.U$$650/B VGND VGND VPWR VPWR
+ final_adder.U$$762/B sky130_fd_sc_hd__and2_1
XTAP_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$661 final_adder.U$$660/B final_adder.U$$557/X final_adder.U$$541/X
+ VGND VGND VPWR VPWR final_adder.U$$661/X sky130_fd_sc_hd__a21o_1
XTAP_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$500 U$$500/A U$$504/B VGND VGND VPWR VPWR U$$500/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$672 final_adder.U$$688/B final_adder.U$$672/B VGND VGND VPWR VPWR
+ final_adder.U$$784/B sky130_fd_sc_hd__and2_1
XU$$511 U$$783/B1 U$$515/A2 U$$650/A1 U$$515/B2 VGND VGND VPWR VPWR U$$512/A sky130_fd_sc_hd__a22o_1
XTAP_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_36_3 dadda_fa_3_36_3/A dadda_fa_3_36_3/B dadda_fa_3_36_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_37_1/B dadda_fa_4_36_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$683 final_adder.U$$682/B final_adder.U$$579/X final_adder.U$$563/X
+ VGND VGND VPWR VPWR final_adder.U$$683/X sky130_fd_sc_hd__a21o_1
XTAP_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$522 U$$522/A U$$528/B VGND VGND VPWR VPWR U$$522/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$694 final_adder.U$$710/B final_adder.U$$694/B VGND VGND VPWR VPWR
+ final_adder.U$$774/A sky130_fd_sc_hd__and2_1
XTAP_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$533 U$$807/A1 U$$537/A2 U$$807/B1 U$$537/B2 VGND VGND VPWR VPWR U$$534/A sky130_fd_sc_hd__a22o_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$544 U$$544/A U$$546/B VGND VGND VPWR VPWR U$$544/X sky130_fd_sc_hd__xor2_1
XU$$555 U$$555/A U$$607/B VGND VGND VPWR VPWR U$$555/X sky130_fd_sc_hd__xor2_1
XTAP_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$566 U$$703/A1 U$$578/A2 U$$20/A1 U$$578/B2 VGND VGND VPWR VPWR U$$567/A sky130_fd_sc_hd__a22o_1
XTAP_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_29_2 dadda_fa_3_29_2/A dadda_fa_3_29_2/B dadda_fa_3_29_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_30_1/A dadda_fa_4_29_2/B sky130_fd_sc_hd__fa_2
XFILLER_17_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$577 U$$577/A U$$579/B VGND VGND VPWR VPWR U$$577/X sky130_fd_sc_hd__xor2_1
XU$$588 U$$997/B1 U$$624/A2 U$$864/A1 U$$624/B2 VGND VGND VPWR VPWR U$$589/A sky130_fd_sc_hd__a22o_1
XFILLER_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$599 U$$599/A U$$617/B VGND VGND VPWR VPWR U$$599/X sky130_fd_sc_hd__xor2_1
XFILLER_60_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1400 U$$2311/B VGND VGND VPWR VPWR U$$2309/B sky130_fd_sc_hd__buf_6
XFILLER_201_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1411 U$$2043/B VGND VGND VPWR VPWR U$$1993/B sky130_fd_sc_hd__buf_6
Xrepeater1422 U$$1832/B VGND VGND VPWR VPWR U$$1840/B sky130_fd_sc_hd__buf_8
XFILLER_153_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1433 U$$1751/B VGND VGND VPWR VPWR U$$1707/B sky130_fd_sc_hd__buf_6
XFILLER_207_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1444 U$$1644/A VGND VGND VPWR VPWR U$$1608/B sky130_fd_sc_hd__buf_8
XFILLER_126_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1455 input14/X VGND VGND VPWR VPWR U$$1507/A sky130_fd_sc_hd__buf_6
XFILLER_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1466 U$$709/A1 VGND VGND VPWR VPWR U$$983/A1 sky130_fd_sc_hd__buf_4
XFILLER_181_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1477 U$$4406/A1 VGND VGND VPWR VPWR U$$4269/A1 sky130_fd_sc_hd__buf_6
XFILLER_154_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1488 input125/X VGND VGND VPWR VPWR U$$431/A1 sky130_fd_sc_hd__buf_4
XFILLER_158_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1499 U$$2324/A1 VGND VGND VPWR VPWR U$$954/A1 sky130_fd_sc_hd__buf_6
XFILLER_41_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_31_2 U$$867/X U$$1000/X U$$1133/X VGND VGND VPWR VPWR dadda_fa_3_32_1/B
+ dadda_fa_3_31_3/B sky130_fd_sc_hd__fa_1
XFILLER_208_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1250 U$$1250/A U$$1270/B VGND VGND VPWR VPWR U$$1250/X sky130_fd_sc_hd__xor2_1
XFILLER_189_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1261 U$$2220/A1 U$$1289/A2 U$$989/A1 U$$1281/B2 VGND VGND VPWR VPWR U$$1262/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1272 U$$1272/A U$$1272/B VGND VGND VPWR VPWR U$$1272/X sky130_fd_sc_hd__xor2_1
XFILLER_189_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1283 U$$461/A1 U$$1289/A2 U$$461/B1 U$$1291/B2 VGND VGND VPWR VPWR U$$1284/A sky130_fd_sc_hd__a22o_1
XFILLER_176_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1294 U$$1294/A U$$1330/B VGND VGND VPWR VPWR U$$1294/X sky130_fd_sc_hd__xor2_1
XFILLER_31_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_5 U$$3365/X U$$3498/X U$$3631/X VGND VGND VPWR VPWR dadda_fa_2_84_3/B
+ dadda_fa_2_83_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_76_4 U$$3085/X U$$3218/X U$$3351/X VGND VGND VPWR VPWR dadda_fa_2_77_1/CIN
+ dadda_fa_2_76_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_502 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_3 U$$3603/X U$$3736/X U$$3869/X VGND VGND VPWR VPWR dadda_fa_2_70_1/B
+ dadda_fa_2_69_4/B sky130_fd_sc_hd__fa_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_46_2 dadda_fa_4_46_2/A dadda_fa_4_46_2/B dadda_fa_4_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_47_0/CIN dadda_fa_5_46_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_39_1 dadda_fa_4_39_1/A dadda_fa_4_39_1/B dadda_fa_4_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/B dadda_fa_5_39_1/B sky130_fd_sc_hd__fa_1
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _200_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_7_16_0 dadda_fa_7_16_0/A dadda_fa_7_16_0/B dadda_fa_7_16_0/CIN VGND VGND
+ VPWR VPWR _313_/D _184_/D sky130_fd_sc_hd__fa_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_239 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_290_ _419_/CLK _290_/D VGND VGND VPWR VPWR _290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_0_58_3 U$$1320/X U$$1453/X VGND VGND VPWR VPWR dadda_fa_1_59_7/CIN dadda_fa_2_58_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_27_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_71_3 U$$1745/X U$$1878/X U$$2011/X VGND VGND VPWR VPWR dadda_fa_1_72_7/CIN
+ dadda_fa_2_71_0/A sky130_fd_sc_hd__fa_1
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_693 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_64_2 U$$933/X U$$1066/X U$$1199/X VGND VGND VPWR VPWR dadda_fa_1_65_6/A
+ dadda_fa_1_64_8/A sky130_fd_sc_hd__fa_1
XTAP_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1056 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_41_1 dadda_fa_3_41_1/A dadda_fa_3_41_1/B dadda_fa_3_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_0/CIN dadda_fa_4_41_2/A sky130_fd_sc_hd__fa_1
XTAP_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_57_1 U$$520/X U$$653/X U$$786/X VGND VGND VPWR VPWR dadda_fa_1_58_7/B
+ dadda_fa_1_57_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$480 final_adder.U$$484/B final_adder.U$$480/B VGND VGND VPWR VPWR
+ final_adder.U$$604/B sky130_fd_sc_hd__and2_1
XTAP_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_34_0 dadda_fa_3_34_0/A dadda_fa_3_34_0/B dadda_fa_3_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_0/B dadda_fa_4_34_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$491 final_adder.U$$490/B final_adder.U$$369/X final_adder.U$$365/X
+ VGND VGND VPWR VPWR final_adder.U$$491/X sky130_fd_sc_hd__a21o_1
XTAP_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$330 U$$330/A1 U$$350/A2 U$$56/B1 U$$350/B2 VGND VGND VPWR VPWR U$$331/A sky130_fd_sc_hd__a22o_1
XTAP_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$341 U$$341/A U$$367/B VGND VGND VPWR VPWR U$$341/X sky130_fd_sc_hd__xor2_1
XTAP_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$352 U$$763/A1 U$$396/A2 U$$763/B1 U$$396/B2 VGND VGND VPWR VPWR U$$353/A sky130_fd_sc_hd__a22o_1
XTAP_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$363 U$$363/A U$$397/B VGND VGND VPWR VPWR U$$363/X sky130_fd_sc_hd__xor2_1
XFILLER_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$374 U$$920/B1 U$$378/A2 U$$787/A1 U$$378/B2 VGND VGND VPWR VPWR U$$375/A sky130_fd_sc_hd__a22o_1
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$385 U$$385/A U$$395/B VGND VGND VPWR VPWR U$$385/X sky130_fd_sc_hd__xor2_1
XFILLER_17_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$396 U$$807/A1 U$$396/A2 U$$807/B1 U$$396/B2 VGND VGND VPWR VPWR U$$397/A sky130_fd_sc_hd__a22o_1
XFILLER_60_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_93_4 U$$4449/X input249/X dadda_fa_2_93_4/CIN VGND VGND VPWR VPWR dadda_fa_3_94_1/CIN
+ dadda_fa_3_93_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1230 input60/X VGND VGND VPWR VPWR U$$4370/B sky130_fd_sc_hd__buf_6
Xrepeater1241 U$$397/B VGND VGND VPWR VPWR U$$351/B sky130_fd_sc_hd__buf_8
XFILLER_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1252 input55/X VGND VGND VPWR VPWR U$$4100/B sky130_fd_sc_hd__buf_6
XFILLER_181_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_86_3 dadda_fa_2_86_3/A dadda_fa_2_86_3/B dadda_fa_2_86_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_1/B dadda_fa_3_86_3/B sky130_fd_sc_hd__fa_1
Xrepeater1263 U$$3875/B VGND VGND VPWR VPWR U$$3903/B sky130_fd_sc_hd__buf_8
XFILLER_114_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1274 U$$3836/A VGND VGND VPWR VPWR U$$3834/B sky130_fd_sc_hd__buf_6
Xrepeater1285 U$$3609/B VGND VGND VPWR VPWR U$$3613/B sky130_fd_sc_hd__buf_6
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1296 U$$3518/B VGND VGND VPWR VPWR U$$3550/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_79_2 dadda_fa_2_79_2/A dadda_fa_2_79_2/B dadda_fa_2_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/A dadda_fa_3_79_3/A sky130_fd_sc_hd__fa_1
XFILLER_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_56_1 dadda_fa_5_56_1/A dadda_fa_5_56_1/B dadda_fa_5_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_57_0/B dadda_fa_7_56_0/A sky130_fd_sc_hd__fa_1
XFILLER_84_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_49_0 dadda_fa_5_49_0/A dadda_fa_5_49_0/B dadda_fa_5_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_50_0/A dadda_fa_6_49_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_23_0 U$$53/X U$$186/X VGND VGND VPWR VPWR dadda_fa_3_24_3/B dadda_fa_4_23_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_209_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_102_1 U$$3004/X U$$3137/X U$$3270/X VGND VGND VPWR VPWR dadda_fa_3_103_2/B
+ dadda_fa_3_102_3/B sky130_fd_sc_hd__fa_1
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1080 U$$1080/A U$$1095/A VGND VGND VPWR VPWR U$$1080/X sky130_fd_sc_hd__xor2_1
XU$$1091 U$$954/A1 U$$1093/A2 U$$1504/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1092/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_123_0 U$$4109/Y U$$4243/X U$$4376/X VGND VGND VPWR VPWR dadda_fa_6_124_0/A
+ dadda_fa_6_123_0/CIN sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_30_clk _255_/CLK VGND VGND VPWR VPWR _412_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_81_2 U$$2031/X U$$2164/X U$$2297/X VGND VGND VPWR VPWR dadda_fa_2_82_1/CIN
+ dadda_fa_2_81_4/B sky130_fd_sc_hd__fa_1
XFILLER_105_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_74_1 U$$2150/X U$$2283/X U$$2416/X VGND VGND VPWR VPWR dadda_fa_2_75_0/CIN
+ dadda_fa_2_74_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_51_0 dadda_fa_4_51_0/A dadda_fa_4_51_0/B dadda_fa_4_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/A dadda_fa_5_51_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_67_0 U$$2535/X U$$2668/X U$$2801/X VGND VGND VPWR VPWR dadda_fa_2_68_0/B
+ dadda_fa_2_67_3/B sky130_fd_sc_hd__fa_1
XFILLER_59_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2709 U$$2709/A1 U$$2607/X U$$2709/B1 U$$2608/X VGND VGND VPWR VPWR U$$2710/A sky130_fd_sc_hd__a22o_1
XFILLER_74_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1055 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_411_ _411_/CLK _411_/D VGND VGND VPWR VPWR _411_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_342_ _342_/CLK _342_/D VGND VGND VPWR VPWR _342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_273_ _401_/CLK _273_/D VGND VGND VPWR VPWR _273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_clk _380_/CLK VGND VGND VPWR VPWR _399_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_96_2 dadda_fa_3_96_2/A dadda_fa_3_96_2/B dadda_fa_3_96_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_1/A dadda_fa_4_96_2/B sky130_fd_sc_hd__fa_1
XFILLER_108_551 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_89_1 dadda_fa_3_89_1/A dadda_fa_3_89_1/B dadda_fa_3_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_0/CIN dadda_fa_4_89_2/A sky130_fd_sc_hd__fa_1
XFILLER_185_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_66_0 dadda_fa_6_66_0/A dadda_fa_6_66_0/B dadda_fa_6_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_67_0/B dadda_fa_7_66_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater908 U$$3648/B1 VGND VGND VPWR VPWR U$$3376/A1 sky130_fd_sc_hd__buf_6
XFILLER_89_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater919 U$$3922/A1 VGND VGND VPWR VPWR U$$84/B1 sky130_fd_sc_hd__buf_6
XFILLER_77_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3696_1752 VGND VGND VPWR VPWR U$$3696_1752/HI U$$3696/B1 sky130_fd_sc_hd__conb_1
XU$$3900 U$$4309/B1 U$$3902/A2 U$$4176/A1 U$$3902/B2 VGND VGND VPWR VPWR U$$3901/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3911 U$$3911/A U$$3971/B VGND VGND VPWR VPWR U$$3911/X sky130_fd_sc_hd__xor2_1
XTAP_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_118_1 U$$4100/X U$$4233/X U$$4366/X VGND VGND VPWR VPWR dadda_fa_5_119_0/CIN
+ dadda_fa_5_118_1/B sky130_fd_sc_hd__fa_1
XFILLER_64_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3922 U$$3922/A1 U$$3926/A2 U$$3922/B1 U$$3926/B2 VGND VGND VPWR VPWR U$$3923/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3933 U$$3933/A U$$3947/B VGND VGND VPWR VPWR U$$3933/X sky130_fd_sc_hd__xor2_1
XFILLER_18_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3944 U$$3944/A1 U$$3946/A2 U$$3944/B1 U$$3946/B2 VGND VGND VPWR VPWR U$$3945/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3955 U$$3955/A U$$3972/A VGND VGND VPWR VPWR U$$3955/X sky130_fd_sc_hd__xor2_1
XTAP_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3966 U$$4375/B1 U$$3966/A2 U$$4103/B1 U$$3966/B2 VGND VGND VPWR VPWR U$$3967/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3977 U$$3975/Y input54/X input53/X U$$3976/X U$$3973/Y VGND VGND VPWR VPWR U$$3977/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_206_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$160 U$$160/A U$$160/B VGND VGND VPWR VPWR U$$160/X sky130_fd_sc_hd__xor2_1
XU$$3988 U$$3988/A U$$4012/B VGND VGND VPWR VPWR U$$3988/X sky130_fd_sc_hd__xor2_1
XTAP_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3999 U$$4273/A1 U$$4035/A2 U$$4273/B1 U$$4035/B2 VGND VGND VPWR VPWR U$$4000/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$171 U$$34/A1 U$$175/A2 U$$36/A1 U$$175/B2 VGND VGND VPWR VPWR U$$172/A sky130_fd_sc_hd__a22o_1
XU$$182 U$$182/A U$$184/B VGND VGND VPWR VPWR U$$182/X sky130_fd_sc_hd__xor2_1
XFILLER_206_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$193 U$$328/B1 U$$217/A2 U$$58/A1 U$$217/B2 VGND VGND VPWR VPWR U$$194/A sky130_fd_sc_hd__a22o_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_12_clk _227_/CLK VGND VGND VPWR VPWR _359_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_91_1 U$$3514/X U$$3647/X U$$3780/X VGND VGND VPWR VPWR dadda_fa_3_92_0/CIN
+ dadda_fa_3_91_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_12_1174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_84_0 U$$4032/X U$$4165/X U$$4298/X VGND VGND VPWR VPWR dadda_fa_3_85_0/B
+ dadda_fa_3_84_2/B sky130_fd_sc_hd__fa_1
Xrepeater1060 U$$3344/A1 VGND VGND VPWR VPWR U$$741/A1 sky130_fd_sc_hd__buf_8
XFILLER_99_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput257 output257/A VGND VGND VPWR VPWR o[0] sky130_fd_sc_hd__buf_2
XFILLER_47_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1071 U$$4027/A1 VGND VGND VPWR VPWR U$$4162/B1 sky130_fd_sc_hd__buf_8
Xoutput268 output268/A VGND VGND VPWR VPWR o[10] sky130_fd_sc_hd__buf_2
Xrepeater1082 U$$50/A1 VGND VGND VPWR VPWR U$$48/B1 sky130_fd_sc_hd__buf_4
Xoutput279 output279/A VGND VGND VPWR VPWR o[11] sky130_fd_sc_hd__buf_2
XFILLER_173_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1093 U$$3747/A1 VGND VGND VPWR VPWR U$$733/A1 sky130_fd_sc_hd__buf_6
XFILLER_114_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_60_7 dadda_fa_1_60_7/A dadda_fa_1_60_7/B dadda_fa_1_60_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_61_2/CIN dadda_fa_2_60_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_6 U$$2773/X U$$2906/X U$$3039/X VGND VGND VPWR VPWR dadda_fa_2_54_2/B
+ dadda_fa_2_53_5/B sky130_fd_sc_hd__fa_1
XFILLER_68_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_46_5 U$$2094/X U$$2227/X U$$2360/X VGND VGND VPWR VPWR dadda_fa_2_47_3/B
+ dadda_fa_2_46_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_70_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_5_0 dadda_fa_7_5_0/A dadda_fa_7_5_0/B dadda_fa_7_5_0/CIN VGND VGND VPWR
+ VPWR _302_/D _173_/D sky130_fd_sc_hd__fa_1
XFILLER_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1109 final_adder.U$$170/B final_adder.U$$941/X VGND VGND VPWR VPWR
+ output368/A sky130_fd_sc_hd__xor2_1
XFILLER_177_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_83_0 dadda_fa_7_83_0/A dadda_fa_7_83_0/B dadda_fa_7_83_0/CIN VGND VGND
+ VPWR VPWR _380_/D _251_/D sky130_fd_sc_hd__fa_2
XFILLER_109_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_99_0 dadda_fa_4_99_0/A dadda_fa_4_99_0/B dadda_fa_4_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/A dadda_fa_5_99_1/A sky130_fd_sc_hd__fa_1
XFILLER_192_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3207 U$$741/A1 U$$3207/A2 U$$3207/B1 U$$3207/B2 VGND VGND VPWR VPWR U$$3208/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1252 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3218 U$$3218/A U$$3256/B VGND VGND VPWR VPWR U$$3218/X sky130_fd_sc_hd__xor2_1
XFILLER_115_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3229 U$$3775/B1 U$$3229/A2 U$$3642/A1 U$$3156/X VGND VGND VPWR VPWR U$$3230/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2506 U$$38/B1 U$$2596/A2 U$$4013/B1 U$$2596/B2 VGND VGND VPWR VPWR U$$2507/A sky130_fd_sc_hd__a22o_1
XFILLER_62_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2517 U$$2517/A U$$2543/B VGND VGND VPWR VPWR U$$2517/X sky130_fd_sc_hd__xor2_1
XU$$2528 U$$3211/B1 U$$2558/A2 U$$3352/A1 U$$2558/B2 VGND VGND VPWR VPWR U$$2529/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2539 U$$2539/A U$$2569/B VGND VGND VPWR VPWR U$$2539/X sky130_fd_sc_hd__xor2_1
XFILLER_64_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1805 U$$709/A1 U$$1839/A2 U$$983/B1 U$$1839/B2 VGND VGND VPWR VPWR U$$1806/A sky130_fd_sc_hd__a22o_1
XU$$1816 U$$1816/A U$$1820/B VGND VGND VPWR VPWR U$$1816/X sky130_fd_sc_hd__xor2_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1827 U$$731/A1 U$$1877/A2 U$$594/B1 U$$1877/B2 VGND VGND VPWR VPWR U$$1828/A sky130_fd_sc_hd__a22o_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1838 U$$1838/A U$$1840/B VGND VGND VPWR VPWR U$$1838/X sky130_fd_sc_hd__xor2_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1849 U$$4452/A1 U$$1915/A2 U$$4454/A1 U$$1915/B2 VGND VGND VPWR VPWR U$$1850/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ _325_/CLK _325_/D VGND VGND VPWR VPWR _325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_579 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_256_ _390_/CLK _256_/D VGND VGND VPWR VPWR _256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_187_ _326_/CLK _187_/D VGND VGND VPWR VPWR _187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_63_5 dadda_fa_2_63_5/A dadda_fa_2_63_5/B dadda_fa_2_63_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_2/A dadda_fa_4_63_0/A sky130_fd_sc_hd__fa_2
XFILLER_85_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater705 U$$3841/X VGND VGND VPWR VPWR U$$3970/B2 sky130_fd_sc_hd__buf_6
XFILLER_1_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater716 U$$3704/X VGND VGND VPWR VPWR U$$3773/B2 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_1_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _208_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater727 U$$3479/B2 VGND VGND VPWR VPWR U$$3453/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_56_4 dadda_fa_2_56_4/A dadda_fa_2_56_4/B dadda_fa_2_56_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_1/CIN dadda_fa_3_56_3/CIN sky130_fd_sc_hd__fa_2
Xrepeater738 U$$3390/B2 VGND VGND VPWR VPWR U$$3416/B2 sky130_fd_sc_hd__buf_6
XU$$4420 U$$4420/A1 U$$4388/X U$$4422/A1 U$$4426/B2 VGND VGND VPWR VPWR U$$4421/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater749 U$$3156/X VGND VGND VPWR VPWR U$$3255/B2 sky130_fd_sc_hd__buf_4
XU$$4431 U$$4431/A U$$4431/B VGND VGND VPWR VPWR U$$4431/X sky130_fd_sc_hd__xor2_1
XU$$4442 U$$4442/A1 U$$4388/X U$$4442/B1 U$$4512/B2 VGND VGND VPWR VPWR U$$4443/A
+ sky130_fd_sc_hd__a22o_1
XU$$4453 U$$4453/A U$$4453/B VGND VGND VPWR VPWR U$$4453/X sky130_fd_sc_hd__xor2_1
XU$$4464 U$$4464/A1 U$$4388/X U$$4466/A1 U$$4476/B2 VGND VGND VPWR VPWR U$$4465/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_49_3 dadda_fa_2_49_3/A dadda_fa_2_49_3/B dadda_fa_2_49_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/B dadda_fa_3_49_3/B sky130_fd_sc_hd__fa_1
XU$$4475 U$$4475/A U$$4475/B VGND VGND VPWR VPWR U$$4475/X sky130_fd_sc_hd__xor2_1
XU$$3730 U$$3730/A U$$3774/B VGND VGND VPWR VPWR U$$3730/X sky130_fd_sc_hd__xor2_1
XFILLER_77_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4486 input106/X U$$4388/X U$$4488/A1 U$$4486/B2 VGND VGND VPWR VPWR U$$4487/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3741 U$$3876/B1 U$$3777/A2 U$$3878/B1 U$$3777/B2 VGND VGND VPWR VPWR U$$3742/A
+ sky130_fd_sc_hd__a22o_1
XU$$4497 U$$4497/A U$$4497/B VGND VGND VPWR VPWR U$$4497/X sky130_fd_sc_hd__xor2_1
XU$$3752 U$$3752/A U$$3754/B VGND VGND VPWR VPWR U$$3752/X sky130_fd_sc_hd__xor2_1
XU$$3763 U$$4309/B1 U$$3773/A2 U$$4176/A1 U$$3773/B2 VGND VGND VPWR VPWR U$$3764/A
+ sky130_fd_sc_hd__a22o_1
XU$$3774 U$$3774/A U$$3774/B VGND VGND VPWR VPWR U$$3774/X sky130_fd_sc_hd__xor2_1
XU$$3785 U$$4333/A1 U$$3813/A2 U$$4333/B1 U$$3813/B2 VGND VGND VPWR VPWR U$$3786/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_19_1 dadda_fa_5_19_1/A dadda_fa_5_19_1/B dadda_fa_5_19_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_20_0/B dadda_fa_7_19_0/A sky130_fd_sc_hd__fa_1
XU$$3796 U$$3796/A U$$3814/B VGND VGND VPWR VPWR U$$3796/X sky130_fd_sc_hd__xor2_1
XFILLER_79_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_51_3 U$$1306/X U$$1439/X U$$1572/X VGND VGND VPWR VPWR dadda_fa_2_52_1/B
+ dadda_fa_2_51_4/B sky130_fd_sc_hd__fa_1
XFILLER_56_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$907 U$$907/A U$$919/B VGND VGND VPWR VPWR U$$907/X sky130_fd_sc_hd__xor2_1
XU$$918 U$$918/A1 U$$918/A2 U$$920/A1 U$$918/B2 VGND VGND VPWR VPWR U$$919/A sky130_fd_sc_hd__a22o_1
XFILLER_16_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_44_2 U$$893/X U$$1026/X U$$1159/X VGND VGND VPWR VPWR dadda_fa_2_45_3/A
+ dadda_fa_2_44_5/A sky130_fd_sc_hd__fa_1
XU$$929 U$$929/A U$$929/B VGND VGND VPWR VPWR U$$929/X sky130_fd_sc_hd__xor2_1
XFILLER_3_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_21_1 dadda_fa_4_21_1/A dadda_fa_4_21_1/B dadda_fa_4_21_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_22_0/B dadda_fa_5_21_1/B sky130_fd_sc_hd__fa_1
XFILLER_71_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_14_0 U$$301/X U$$434/X U$$567/X VGND VGND VPWR VPWR dadda_fa_5_15_0/A
+ dadda_fa_5_14_1/A sky130_fd_sc_hd__fa_1
XFILLER_169_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_78_0_1871 VGND VGND VPWR VPWR dadda_ha_0_78_0/A dadda_ha_0_78_0_1871/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4489_1821 VGND VGND VPWR VPWR U$$4489_1821/HI U$$4489/B sky130_fd_sc_hd__conb_1
Xdadda_fa_3_66_3 dadda_fa_3_66_3/A dadda_fa_3_66_3/B dadda_fa_3_66_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_67_1/B dadda_fa_4_66_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_59_2 dadda_fa_3_59_2/A dadda_fa_3_59_2/B dadda_fa_3_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_1/A dadda_fa_4_59_2/B sky130_fd_sc_hd__fa_1
XFILLER_120_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3004 U$$3004/A U$$3013/A VGND VGND VPWR VPWR U$$3004/X sky130_fd_sc_hd__xor2_1
XU$$3015 input39/X VGND VGND VPWR VPWR U$$3017/B sky130_fd_sc_hd__inv_1
XFILLER_75_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_29_0 dadda_fa_6_29_0/A dadda_fa_6_29_0/B dadda_fa_6_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_30_0/B dadda_fa_7_29_0/CIN sky130_fd_sc_hd__fa_1
XU$$3026 U$$3026/A1 U$$3060/A2 U$$3028/A1 U$$3060/B2 VGND VGND VPWR VPWR U$$3027/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3037 U$$3037/A U$$3125/B VGND VGND VPWR VPWR U$$3037/X sky130_fd_sc_hd__xor2_1
XFILLER_35_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2303 U$$2303/A U$$2303/B VGND VGND VPWR VPWR U$$2303/X sky130_fd_sc_hd__xor2_1
XU$$3048 U$$4144/A1 U$$3082/A2 U$$4144/B1 U$$3082/B2 VGND VGND VPWR VPWR U$$3049/A
+ sky130_fd_sc_hd__a22o_1
XU$$2314 U$$4506/A1 U$$2316/A2 U$$4369/B1 U$$2316/B2 VGND VGND VPWR VPWR U$$2315/A
+ sky130_fd_sc_hd__a22o_1
XU$$3059 U$$3059/A U$$3077/B VGND VGND VPWR VPWR U$$3059/X sky130_fd_sc_hd__xor2_1
XU$$2325 U$$2325/A U$$2328/A VGND VGND VPWR VPWR U$$2325/X sky130_fd_sc_hd__xor2_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2336 U$$2336/A U$$2366/B VGND VGND VPWR VPWR U$$2336/X sky130_fd_sc_hd__xor2_1
XU$$1602 U$$1602/A U$$1608/B VGND VGND VPWR VPWR U$$1602/X sky130_fd_sc_hd__xor2_1
XU$$2347 U$$2621/A1 U$$2359/A2 U$$2623/A1 U$$2359/B2 VGND VGND VPWR VPWR U$$2348/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2358 U$$2358/A U$$2360/B VGND VGND VPWR VPWR U$$2358/X sky130_fd_sc_hd__xor2_1
XU$$1613 U$$2159/B1 U$$1635/A2 U$$2026/A1 U$$1635/B2 VGND VGND VPWR VPWR U$$1614/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2369 U$$38/B1 U$$2463/A2 U$$179/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2370/A sky130_fd_sc_hd__a22o_1
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1624 U$$1624/A U$$1628/B VGND VGND VPWR VPWR U$$1624/X sky130_fd_sc_hd__xor2_1
XU$$1635 U$$2044/B1 U$$1635/A2 U$$950/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1636/A
+ sky130_fd_sc_hd__a22o_1
XU$$1646 U$$1779/B VGND VGND VPWR VPWR U$$1646/Y sky130_fd_sc_hd__inv_1
XFILLER_91_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1657 U$$1657/A U$$1689/B VGND VGND VPWR VPWR U$$1657/X sky130_fd_sc_hd__xor2_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1668 U$$983/A1 U$$1706/A2 U$$983/B1 U$$1706/B2 VGND VGND VPWR VPWR U$$1669/A sky130_fd_sc_hd__a22o_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1679 U$$1679/A U$$1679/B VGND VGND VPWR VPWR U$$1679/X sky130_fd_sc_hd__xor2_1
XFILLER_202_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_308_ _314_/CLK _308_/D VGND VGND VPWR VPWR _308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_239_ _239_/CLK _239_/D VGND VGND VPWR VPWR _239_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_200_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_61_2 dadda_fa_2_61_2/A dadda_fa_2_61_2/B dadda_fa_2_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/A dadda_fa_3_61_3/A sky130_fd_sc_hd__fa_1
XFILLER_170_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater502 U$$3155/X VGND VGND VPWR VPWR U$$3229/A2 sky130_fd_sc_hd__buf_6
XFILLER_97_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$309 final_adder.U$$308/B final_adder.U$$183/X final_adder.U$$181/X
+ VGND VGND VPWR VPWR final_adder.U$$309/X sky130_fd_sc_hd__a21o_1
Xrepeater513 U$$2949/A2 VGND VGND VPWR VPWR U$$2921/A2 sky130_fd_sc_hd__buf_4
Xrepeater524 U$$394/A2 VGND VGND VPWR VPWR U$$366/A2 sky130_fd_sc_hd__buf_6
XFILLER_66_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_54_1 dadda_fa_2_54_1/A dadda_fa_2_54_1/B dadda_fa_2_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_0/CIN dadda_fa_3_54_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater535 U$$2744/X VGND VGND VPWR VPWR U$$2844/A2 sky130_fd_sc_hd__buf_6
Xrepeater546 U$$2470/X VGND VGND VPWR VPWR U$$2588/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_211_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater557 U$$2449/A2 VGND VGND VPWR VPWR U$$2459/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_66_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater568 U$$2169/A2 VGND VGND VPWR VPWR U$$2091/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_31_0 dadda_fa_5_31_0/A dadda_fa_5_31_0/B dadda_fa_5_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_32_0/A dadda_fa_6_31_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_47_0 U$$2761/X U$$2894/X U$$3027/X VGND VGND VPWR VPWR dadda_fa_3_48_0/B
+ dadda_fa_3_47_2/B sky130_fd_sc_hd__fa_1
Xrepeater579 U$$2046/A2 VGND VGND VPWR VPWR U$$2022/A2 sky130_fd_sc_hd__buf_6
XU$$4250 input60/X U$$4250/B VGND VGND VPWR VPWR U$$4250/X sky130_fd_sc_hd__and2_1
XU$$4261 U$$4398/A1 U$$4381/A2 U$$4400/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4262/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4272 U$$4272/A U$$4278/B VGND VGND VPWR VPWR U$$4272/X sky130_fd_sc_hd__xor2_1
XU$$4283 input70/X U$$4327/A2 input71/X U$$4327/B2 VGND VGND VPWR VPWR U$$4284/A sky130_fd_sc_hd__a22o_1
XFILLER_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4294 U$$4294/A U$$4294/B VGND VGND VPWR VPWR U$$4294/X sky130_fd_sc_hd__xor2_1
XU$$3560 U$$3560/A U$$3561/A VGND VGND VPWR VPWR U$$3560/X sky130_fd_sc_hd__xor2_1
XFILLER_198_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3571 U$$3571/A U$$3609/B VGND VGND VPWR VPWR U$$3571/X sky130_fd_sc_hd__xor2_1
XFILLER_53_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3582 U$$4404/A1 U$$3612/A2 U$$4406/A1 U$$3612/B2 VGND VGND VPWR VPWR U$$3583/A
+ sky130_fd_sc_hd__a22o_1
XU$$3593 U$$3593/A U$$3613/B VGND VGND VPWR VPWR U$$3593/X sky130_fd_sc_hd__xor2_1
XFILLER_41_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2870 input122/X U$$2874/A2 U$$3555/B1 U$$2874/B2 VGND VGND VPWR VPWR U$$2871/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_8_1 U$$579/B input245/X dadda_ha_4_8_0/SUM VGND VGND VPWR VPWR dadda_fa_6_9_0/B
+ dadda_fa_7_8_0/A sky130_fd_sc_hd__fa_1
XFILLER_80_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2881 U$$2879/Y input37/X input36/X U$$2880/X U$$2877/Y VGND VGND VPWR VPWR U$$2881/X
+ sky130_fd_sc_hd__a32o_1
XU$$2892 U$$2892/A U$$2922/B VGND VGND VPWR VPWR U$$2892/X sky130_fd_sc_hd__xor2_1
XFILLER_21_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1025 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_76_2 dadda_fa_4_76_2/A dadda_fa_4_76_2/B dadda_fa_4_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_77_0/CIN dadda_fa_5_76_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_69_1 dadda_fa_4_69_1/A dadda_fa_4_69_1/B dadda_fa_4_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/B dadda_fa_5_69_1/B sky130_fd_sc_hd__fa_1
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_46_0 dadda_fa_7_46_0/A dadda_fa_7_46_0/B dadda_fa_7_46_0/CIN VGND VGND
+ VPWR VPWR _343_/D _214_/D sky130_fd_sc_hd__fa_2
XTAP_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$821 final_adder.U$$788/A final_adder.U$$621/X final_adder.U$$709/X
+ VGND VGND VPWR VPWR final_adder.U$$821/X sky130_fd_sc_hd__a21o_1
XFILLER_25_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$843 final_adder.U$$746/X final_adder.U$$811/X final_adder.U$$747/X
+ VGND VGND VPWR VPWR final_adder.U$$843/X sky130_fd_sc_hd__a21o_2
XTAP_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$865 final_adder.U$$768/X final_adder.U$$833/X final_adder.U$$769/X
+ VGND VGND VPWR VPWR final_adder.U$$865/X sky130_fd_sc_hd__a21o_2
XU$$704 U$$704/A U$$712/B VGND VGND VPWR VPWR U$$704/X sky130_fd_sc_hd__xor2_1
XFILLER_21_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$715 U$$850/B1 U$$739/A2 U$$717/A1 U$$739/B2 VGND VGND VPWR VPWR U$$716/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$887 final_adder.U$$790/X final_adder.U$$623/X final_adder.U$$791/X
+ VGND VGND VPWR VPWR final_adder.U$$887/X sky130_fd_sc_hd__a21o_1
XU$$726 U$$726/A U$$750/B VGND VGND VPWR VPWR U$$726/X sky130_fd_sc_hd__xor2_1
XFILLER_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$737 U$$52/A1 U$$749/A2 U$$52/B1 U$$749/B2 VGND VGND VPWR VPWR U$$738/A sky130_fd_sc_hd__a22o_1
XU$$748 U$$748/A U$$750/B VGND VGND VPWR VPWR U$$748/X sky130_fd_sc_hd__xor2_1
XFILLER_204_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$759 U$$896/A1 U$$759/A2 U$$759/B1 U$$759/B2 VGND VGND VPWR VPWR U$$760/A sky130_fd_sc_hd__a22o_1
XFILLER_83_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_831 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1604 input111/X VGND VGND VPWR VPWR U$$3944/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA_9 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1615 U$$4492/A1 VGND VGND VPWR VPWR U$$2848/A1 sky130_fd_sc_hd__buf_4
XFILLER_32_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1626 input11/X VGND VGND VPWR VPWR U$$1366/B sky130_fd_sc_hd__buf_8
XFILLER_152_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1637 U$$4077/B1 VGND VGND VPWR VPWR U$$654/A1 sky130_fd_sc_hd__buf_4
XFILLER_180_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1648 U$$2568/B1 VGND VGND VPWR VPWR U$$2842/B1 sky130_fd_sc_hd__buf_6
Xrepeater1659 U$$4484/B1 VGND VGND VPWR VPWR U$$3116/A1 sky130_fd_sc_hd__buf_6
XFILLER_152_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_71_1 dadda_fa_3_71_1/A dadda_fa_3_71_1/B dadda_fa_3_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_0/CIN dadda_fa_4_71_2/A sky130_fd_sc_hd__fa_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_64_0 dadda_fa_3_64_0/A dadda_fa_3_64_0/B dadda_fa_3_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_0/B dadda_fa_4_64_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_1043 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2100 U$$2100/A U$$2100/B VGND VGND VPWR VPWR U$$2100/X sky130_fd_sc_hd__xor2_1
XFILLER_35_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2111 U$$3481/A1 U$$2113/A2 U$$3618/B1 U$$2113/B2 VGND VGND VPWR VPWR U$$2112/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_100_1 dadda_fa_4_100_1/A dadda_fa_4_100_1/B dadda_fa_4_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/B dadda_fa_5_100_1/B sky130_fd_sc_hd__fa_1
XFILLER_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2122 U$$2122/A U$$2150/B VGND VGND VPWR VPWR U$$2122/X sky130_fd_sc_hd__xor2_1
XU$$2133 U$$3366/A1 U$$2177/A2 U$$3366/B1 U$$2177/B2 VGND VGND VPWR VPWR U$$2134/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2144 U$$2144/A U$$2150/B VGND VGND VPWR VPWR U$$2144/X sky130_fd_sc_hd__xor2_1
XFILLER_23_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1410 U$$997/B1 U$$1434/A2 U$$864/A1 U$$1434/B2 VGND VGND VPWR VPWR U$$1411/A sky130_fd_sc_hd__a22o_1
XU$$2155 U$$2701/B1 U$$2189/A2 U$$2292/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2156/A
+ sky130_fd_sc_hd__a22o_1
XU$$1421 U$$1421/A U$$1459/B VGND VGND VPWR VPWR U$$1421/X sky130_fd_sc_hd__xor2_1
XU$$2166 U$$2166/A U$$2184/B VGND VGND VPWR VPWR U$$2166/X sky130_fd_sc_hd__xor2_1
XU$$2177 U$$2312/B1 U$$2177/A2 U$$4508/A1 U$$2177/B2 VGND VGND VPWR VPWR U$$2178/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1432 U$$610/A1 U$$1434/A2 U$$610/B1 U$$1434/B2 VGND VGND VPWR VPWR U$$1433/A sky130_fd_sc_hd__a22o_1
XU$$2188 U$$2188/A U$$2191/A VGND VGND VPWR VPWR U$$2188/X sky130_fd_sc_hd__xor2_1
XU$$1443 U$$1443/A U$$1449/B VGND VGND VPWR VPWR U$$1443/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1454 U$$2550/A1 U$$1462/A2 U$$2415/A1 U$$1462/B2 VGND VGND VPWR VPWR U$$1455/A
+ sky130_fd_sc_hd__a22o_1
XU$$2199 U$$2199/A U$$2227/B VGND VGND VPWR VPWR U$$2199/X sky130_fd_sc_hd__xor2_1
XU$$1465 U$$1465/A U$$1506/A VGND VGND VPWR VPWR U$$1465/X sky130_fd_sc_hd__xor2_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1476 U$$2159/B1 U$$1374/X U$$2026/A1 U$$1375/X VGND VGND VPWR VPWR U$$1477/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_7_121_0 dadda_fa_7_121_0/A dadda_fa_7_121_0/B dadda_fa_7_121_0/CIN VGND
+ VGND VPWR VPWR _418_/D _289_/D sky130_fd_sc_hd__fa_1
XU$$1487 U$$1487/A U$$1501/B VGND VGND VPWR VPWR U$$1487/X sky130_fd_sc_hd__xor2_1
XFILLER_176_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1498 U$$2318/B1 U$$1502/A2 U$$950/B1 U$$1502/B2 VGND VGND VPWR VPWR U$$1499/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_86_1 dadda_fa_5_86_1/A dadda_fa_5_86_1/B dadda_fa_5_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_87_0/B dadda_fa_7_86_0/A sky130_fd_sc_hd__fa_2
XFILLER_117_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_79_0 dadda_fa_5_79_0/A dadda_fa_5_79_0/B dadda_fa_5_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_80_0/A dadda_fa_6_79_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_78_8 U$$4419/X input232/X dadda_fa_1_78_8/CIN VGND VGND VPWR VPWR dadda_fa_2_79_3/A
+ dadda_fa_3_78_0/A sky130_fd_sc_hd__fa_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$106 _402_/Q _274_/Q VGND VGND VPWR VPWR final_adder.U$$919/B1 final_adder.U$$148/A
+ sky130_fd_sc_hd__ha_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$117 _413_/Q _285_/Q VGND VGND VPWR VPWR final_adder.U$$139/B1 final_adder.U$$138/B
+ sky130_fd_sc_hd__ha_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$139 final_adder.U$$138/B final_adder.U$$909/B1 final_adder.U$$139/B1
+ VGND VGND VPWR VPWR final_adder.U$$139/X sky130_fd_sc_hd__a21o_1
XFILLER_39_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater387 U$$1057/A2 VGND VGND VPWR VPWR U$$979/A2 sky130_fd_sc_hd__buf_4
XFILLER_26_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater398 U$$938/A2 VGND VGND VPWR VPWR U$$950/A2 sky130_fd_sc_hd__buf_8
XFILLER_211_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4080 U$$4080/A U$$4080/B VGND VGND VPWR VPWR U$$4080/X sky130_fd_sc_hd__xor2_1
XFILLER_25_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4091 input115/X U$$4101/A2 U$$4504/A1 U$$4101/B2 VGND VGND VPWR VPWR U$$4092/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3390 U$$650/A1 U$$3394/A2 U$$3801/B1 U$$3390/B2 VGND VGND VPWR VPWR U$$3391/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_81_0 dadda_fa_4_81_0/A dadda_fa_4_81_0/B dadda_fa_4_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/A dadda_fa_5_81_1/A sky130_fd_sc_hd__fa_1
XFILLER_107_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_102_3 dadda_fa_3_102_3/A dadda_fa_3_102_3/B dadda_fa_3_102_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_103_1/B dadda_fa_4_102_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_123_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput102 b[43] VGND VGND VPWR VPWR input102/X sky130_fd_sc_hd__buf_6
XFILLER_49_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput113 b[53] VGND VGND VPWR VPWR input113/X sky130_fd_sc_hd__buf_6
XFILLER_114_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput124 b[63] VGND VGND VPWR VPWR input124/X sky130_fd_sc_hd__buf_6
XTAP_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput135 c[105] VGND VGND VPWR VPWR input135/X sky130_fd_sc_hd__buf_4
XFILLER_102_162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput146 c[115] VGND VGND VPWR VPWR input146/X sky130_fd_sc_hd__clkbuf_4
XTAP_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput157 c[125] VGND VGND VPWR VPWR input157/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 c[1] VGND VGND VPWR VPWR input168/X sky130_fd_sc_hd__clkbuf_4
XTAP_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$640 final_adder.U$$656/B final_adder.U$$640/B VGND VGND VPWR VPWR
+ final_adder.U$$752/B sky130_fd_sc_hd__and2_1
XTAP_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 c[2] VGND VGND VPWR VPWR input179/X sky130_fd_sc_hd__clkbuf_4
XFILLER_57_750 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$651 final_adder.U$$650/B final_adder.U$$547/X final_adder.U$$531/X
+ VGND VGND VPWR VPWR final_adder.U$$651/X sky130_fd_sc_hd__a21o_1
XTAP_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$662 final_adder.U$$678/B final_adder.U$$662/B VGND VGND VPWR VPWR
+ final_adder.U$$774/B sky130_fd_sc_hd__and2_1
XTAP_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_109_0 dadda_fa_6_109_0/A dadda_fa_6_109_0/B dadda_fa_6_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_110_0/B dadda_fa_7_109_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$501 U$$773/B1 U$$527/A2 U$$640/A1 U$$527/B2 VGND VGND VPWR VPWR U$$502/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$673 final_adder.U$$672/B final_adder.U$$569/X final_adder.U$$553/X
+ VGND VGND VPWR VPWR final_adder.U$$673/X sky130_fd_sc_hd__a21o_1
XTAP_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$512 U$$512/A U$$516/B VGND VGND VPWR VPWR U$$512/X sky130_fd_sc_hd__xor2_1
XTAP_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$684 final_adder.U$$700/B final_adder.U$$684/B VGND VGND VPWR VPWR
+ final_adder.U$$796/B sky130_fd_sc_hd__and2_1
XTAP_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$523 U$$660/A1 U$$415/X U$$660/B1 U$$416/X VGND VGND VPWR VPWR U$$524/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$695 final_adder.U$$694/B final_adder.U$$591/X final_adder.U$$575/X
+ VGND VGND VPWR VPWR final_adder.U$$695/X sky130_fd_sc_hd__a21o_1
XFILLER_186_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$534 U$$534/A U$$536/B VGND VGND VPWR VPWR U$$534/X sky130_fd_sc_hd__xor2_1
XFILLER_186_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$545 U$$817/B1 U$$415/X U$$545/B1 U$$416/X VGND VGND VPWR VPWR U$$546/A sky130_fd_sc_hd__a22o_1
XU$$556 U$$967/A1 U$$578/A2 U$$969/A1 U$$578/B2 VGND VGND VPWR VPWR U$$557/A sky130_fd_sc_hd__a22o_1
XTAP_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$567 U$$567/A U$$579/B VGND VGND VPWR VPWR U$$567/X sky130_fd_sc_hd__xor2_1
XTAP_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_29_3 dadda_fa_3_29_3/A dadda_fa_3_29_3/B dadda_fa_3_29_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_30_1/B dadda_fa_4_29_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_60_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$578 U$$578/A1 U$$578/A2 U$$717/A1 U$$578/B2 VGND VGND VPWR VPWR U$$579/A sky130_fd_sc_hd__a22o_1
XFILLER_60_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$589 U$$589/A U$$625/B VGND VGND VPWR VPWR U$$589/X sky130_fd_sc_hd__xor2_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_96_0 dadda_fa_6_96_0/A dadda_fa_6_96_0/B dadda_fa_6_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_97_0/B dadda_fa_7_96_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_201_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1401 input27/X VGND VGND VPWR VPWR U$$2311/B sky130_fd_sc_hd__buf_4
Xrepeater1412 input22/X VGND VGND VPWR VPWR U$$2043/B sky130_fd_sc_hd__buf_6
Xrepeater1423 U$$1880/B VGND VGND VPWR VPWR U$$1832/B sky130_fd_sc_hd__buf_12
Xrepeater1434 U$$1751/B VGND VGND VPWR VPWR U$$1721/B sky130_fd_sc_hd__buf_6
XFILLER_114_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1445 U$$1644/A VGND VGND VPWR VPWR U$$1638/B sky130_fd_sc_hd__buf_8
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1456 U$$983/B1 VGND VGND VPWR VPWR U$$985/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1467 U$$3584/B1 VGND VGND VPWR VPWR U$$2625/B1 sky130_fd_sc_hd__clkbuf_4
Xrepeater1478 U$$842/B1 VGND VGND VPWR VPWR U$$22/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_4_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1489 U$$956/A1 VGND VGND VPWR VPWR U$$817/B1 sky130_fd_sc_hd__buf_4
XFILLER_154_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$5_1836 VGND VGND VPWR VPWR U$$5_1836/HI U$$5/A2 sky130_fd_sc_hd__conb_1
Xdadda_ha_2_32_5 U$$2066/X U$$2199/X VGND VGND VPWR VPWR dadda_fa_3_33_2/A dadda_fa_4_32_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_39_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_31_3 U$$1266/X U$$1399/X U$$1532/X VGND VGND VPWR VPWR dadda_fa_3_32_1/CIN
+ dadda_fa_3_31_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1240 U$$1240/A U$$1272/B VGND VGND VPWR VPWR U$$1240/X sky130_fd_sc_hd__xor2_1
XU$$1251 U$$1799/A1 U$$1271/A2 U$$1799/B1 U$$1281/B2 VGND VGND VPWR VPWR U$$1252/A
+ sky130_fd_sc_hd__a22o_1
XU$$1262 U$$1262/A U$$1286/B VGND VGND VPWR VPWR U$$1262/X sky130_fd_sc_hd__xor2_1
XU$$1273 U$$999/A1 U$$1311/A2 U$$179/A1 U$$1307/B2 VGND VGND VPWR VPWR U$$1274/A sky130_fd_sc_hd__a22o_1
XFILLER_206_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1284 U$$1284/A U$$1330/B VGND VGND VPWR VPWR U$$1284/X sky130_fd_sc_hd__xor2_1
XFILLER_148_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1295 U$$2391/A1 U$$1323/A2 U$$3213/B1 U$$1349/B2 VGND VGND VPWR VPWR U$$1296/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_83_6 U$$3764/X U$$3897/X U$$4030/X VGND VGND VPWR VPWR dadda_fa_2_84_3/CIN
+ dadda_fa_3_83_0/A sky130_fd_sc_hd__fa_1
XFILLER_104_438 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_76_5 U$$3484/X U$$3617/X U$$3750/X VGND VGND VPWR VPWR dadda_fa_2_77_2/A
+ dadda_fa_2_76_5/A sky130_fd_sc_hd__fa_1
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_4 U$$4002/X U$$4135/X U$$4268/X VGND VGND VPWR VPWR dadda_fa_2_70_1/CIN
+ dadda_fa_2_69_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_85_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_39_2 dadda_fa_4_39_2/A dadda_fa_4_39_2/B dadda_fa_4_39_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_40_0/CIN dadda_fa_5_39_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_207 _200_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_218 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 _251_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_46 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_414 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1250 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_100_0 U$$4330/X U$$4463/X input130/X VGND VGND VPWR VPWR dadda_fa_4_101_0/B
+ dadda_fa_4_100_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_867 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_64_3 U$$1332/X U$$1465/X U$$1598/X VGND VGND VPWR VPWR dadda_fa_1_65_6/B
+ dadda_fa_1_64_8/B sky130_fd_sc_hd__fa_1
XTAP_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_41_2 dadda_fa_3_41_2/A dadda_fa_3_41_2/B dadda_fa_3_41_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_1/A dadda_fa_4_41_2/B sky130_fd_sc_hd__fa_1
XFILLER_76_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$470 final_adder.U$$474/B final_adder.U$$470/B VGND VGND VPWR VPWR
+ final_adder.U$$594/B sky130_fd_sc_hd__and2_1
XTAP_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$481 final_adder.U$$480/B final_adder.U$$359/X final_adder.U$$355/X
+ VGND VGND VPWR VPWR final_adder.U$$481/X sky130_fd_sc_hd__a21o_1
XTAP_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$320 U$$731/A1 U$$350/A2 U$$733/A1 U$$350/B2 VGND VGND VPWR VPWR U$$321/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_34_1 dadda_fa_3_34_1/A dadda_fa_3_34_1/B dadda_fa_3_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_0/CIN dadda_fa_4_34_2/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$492 final_adder.U$$496/B final_adder.U$$492/B VGND VGND VPWR VPWR
+ final_adder.U$$616/B sky130_fd_sc_hd__and2_1
XTAP_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$331 U$$331/A U$$351/B VGND VGND VPWR VPWR U$$331/X sky130_fd_sc_hd__xor2_1
XTAP_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$342 U$$342/A1 U$$366/A2 U$$70/A1 U$$366/B2 VGND VGND VPWR VPWR U$$343/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_11_0 dadda_fa_6_11_0/A dadda_fa_6_11_0/B dadda_fa_6_11_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_12_0/B dadda_fa_7_11_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$353 U$$353/A U$$397/B VGND VGND VPWR VPWR U$$353/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_27_0 U$$1125/X U$$1258/X U$$1391/X VGND VGND VPWR VPWR dadda_fa_4_28_0/B
+ dadda_fa_4_27_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$364 U$$90/A1 U$$396/A2 U$$92/A1 U$$396/B2 VGND VGND VPWR VPWR U$$365/A sky130_fd_sc_hd__a22o_1
XFILLER_199_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$375 U$$375/A U$$377/B VGND VGND VPWR VPWR U$$375/X sky130_fd_sc_hd__xor2_1
XU$$386 U$$521/B1 U$$394/A2 U$$660/B1 U$$394/B2 VGND VGND VPWR VPWR U$$387/A sky130_fd_sc_hd__a22o_1
XU$$397 U$$397/A U$$397/B VGND VGND VPWR VPWR U$$397/X sky130_fd_sc_hd__xor2_1
XFILLER_199_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_93_5 dadda_fa_2_93_5/A dadda_fa_2_93_5/B dadda_fa_2_93_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_94_2/A dadda_fa_4_93_0/A sky130_fd_sc_hd__fa_1
Xrepeater1220 U$$528/B VGND VGND VPWR VPWR U$$504/B sky130_fd_sc_hd__buf_8
Xrepeater1231 input60/X VGND VGND VPWR VPWR U$$4382/B sky130_fd_sc_hd__buf_8
XFILLER_141_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1242 U$$411/A VGND VGND VPWR VPWR U$$397/B sky130_fd_sc_hd__buf_6
Xrepeater1253 U$$4044/B VGND VGND VPWR VPWR U$$4012/B sky130_fd_sc_hd__buf_6
XFILLER_153_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1264 U$$3909/B VGND VGND VPWR VPWR U$$3875/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_86_4 dadda_fa_2_86_4/A dadda_fa_2_86_4/B dadda_fa_2_86_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_1/CIN dadda_fa_3_86_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1275 input51/X VGND VGND VPWR VPWR U$$3836/A sky130_fd_sc_hd__buf_4
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1286 U$$3697/B VGND VGND VPWR VPWR U$$3609/B sky130_fd_sc_hd__buf_6
Xrepeater1297 U$$3518/B VGND VGND VPWR VPWR U$$3561/A sky130_fd_sc_hd__buf_8
XU$$2198_1729 VGND VGND VPWR VPWR U$$2198_1729/HI U$$2198/A1 sky130_fd_sc_hd__conb_1
Xdadda_fa_2_79_3 dadda_fa_2_79_3/A dadda_fa_2_79_3/B dadda_fa_2_79_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/B dadda_fa_3_79_3/B sky130_fd_sc_hd__fa_1
XFILLER_45_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_49_1 dadda_fa_5_49_1/A dadda_fa_5_49_1/B dadda_fa_5_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_50_0/B dadda_fa_7_49_0/A sky130_fd_sc_hd__fa_1
XFILLER_80_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_102_2 U$$3403/X U$$3536/X U$$3669/X VGND VGND VPWR VPWR dadda_fa_3_103_2/CIN
+ dadda_fa_3_102_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_208_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_92_0_1858 VGND VGND VPWR VPWR dadda_fa_1_92_0/A dadda_fa_1_92_0_1858/LO
+ sky130_fd_sc_hd__conb_1
XU$$1070 U$$1070/A U$$962/A VGND VGND VPWR VPWR U$$1070/X sky130_fd_sc_hd__xor2_1
XFILLER_143_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1081 U$$1764/B1 U$$1093/A2 U$$946/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1082/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1092 U$$1092/A U$$1095/A VGND VGND VPWR VPWR U$$1092/X sky130_fd_sc_hd__xor2_1
XFILLER_148_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_123_1 U$$4509/X input155/X dadda_fa_5_123_1/CIN VGND VGND VPWR VPWR dadda_fa_6_124_0/B
+ dadda_fa_7_123_0/A sky130_fd_sc_hd__fa_1
XFILLER_13_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_116_0 dadda_fa_5_116_0/A dadda_fa_5_116_0/B dadda_fa_5_116_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_117_0/A dadda_fa_6_116_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_81_3 U$$2430/X U$$2563/X U$$2696/X VGND VGND VPWR VPWR dadda_fa_2_82_2/A
+ dadda_fa_2_81_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_137_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_74_2 U$$2549/X U$$2682/X U$$2815/X VGND VGND VPWR VPWR dadda_fa_2_75_1/A
+ dadda_fa_2_74_4/A sky130_fd_sc_hd__fa_1
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_51_1 dadda_fa_4_51_1/A dadda_fa_4_51_1/B dadda_fa_4_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/B dadda_fa_5_51_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_67_1 U$$2934/X U$$3067/X U$$3200/X VGND VGND VPWR VPWR dadda_fa_2_68_0/CIN
+ dadda_fa_2_67_3/CIN sky130_fd_sc_hd__fa_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_44_0 dadda_fa_4_44_0/A dadda_fa_4_44_0/B dadda_fa_4_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/A dadda_fa_5_44_1/A sky130_fd_sc_hd__fa_1
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_303 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1067 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ _411_/CLK _410_/D VGND VGND VPWR VPWR _410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_341_ _342_/CLK _341_/D VGND VGND VPWR VPWR _341_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_272_ _401_/CLK _272_/D VGND VGND VPWR VPWR _272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_96_3 dadda_fa_3_96_3/A dadda_fa_3_96_3/B dadda_fa_3_96_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_97_1/B dadda_fa_4_96_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_6_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_89_2 dadda_fa_3_89_2/A dadda_fa_3_89_2/B dadda_fa_3_89_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_1/A dadda_fa_4_89_2/B sky130_fd_sc_hd__fa_1
XFILLER_163_691 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_706 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_59_0 dadda_fa_6_59_0/A dadda_fa_6_59_0/B dadda_fa_6_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_60_0/B dadda_fa_7_59_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater909 U$$4333/B1 VGND VGND VPWR VPWR U$$3648/B1 sky130_fd_sc_hd__buf_6
XFILLER_110_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_62_0 U$$131/X U$$264/X U$$397/X VGND VGND VPWR VPWR dadda_fa_1_63_5/B
+ dadda_fa_1_62_7/B sky130_fd_sc_hd__fa_1
XU$$3901 U$$3901/A U$$3903/B VGND VGND VPWR VPWR U$$3901/X sky130_fd_sc_hd__xor2_1
XFILLER_76_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3912 input92/X U$$3966/A2 U$$4049/B1 U$$3966/B2 VGND VGND VPWR VPWR U$$3913/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3923 U$$3923/A U$$3927/B VGND VGND VPWR VPWR U$$3923/X sky130_fd_sc_hd__xor2_1
XU$$3934 U$$4343/B1 U$$3946/A2 U$$4210/A1 U$$3946/B2 VGND VGND VPWR VPWR U$$3935/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3945 U$$3945/A U$$3947/B VGND VGND VPWR VPWR U$$3945/X sky130_fd_sc_hd__xor2_1
XTAP_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3956 U$$4504/A1 U$$3968/A2 U$$4095/A1 U$$3968/B2 VGND VGND VPWR VPWR U$$3957/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3967 U$$3967/A U$$3967/B VGND VGND VPWR VPWR U$$3967/X sky130_fd_sc_hd__xor2_1
XFILLER_166_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3978 U$$3976/B input53/X input54/X U$$3973/Y VGND VGND VPWR VPWR U$$3978/X sky130_fd_sc_hd__a22o_2
XU$$150 U$$150/A U$$160/B VGND VGND VPWR VPWR U$$150/X sky130_fd_sc_hd__xor2_1
XTAP_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3989 U$$4400/A1 U$$4011/A2 U$$4402/A1 U$$4011/B2 VGND VGND VPWR VPWR U$$3990/A
+ sky130_fd_sc_hd__a22o_1
XU$$161 U$$24/A1 U$$175/A2 U$$26/A1 U$$175/B2 VGND VGND VPWR VPWR U$$162/A sky130_fd_sc_hd__a22o_1
XTAP_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$172 U$$172/A U$$176/B VGND VGND VPWR VPWR U$$172/X sky130_fd_sc_hd__xor2_1
XFILLER_60_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$183 U$$46/A1 U$$209/A2 U$$48/A1 U$$209/B2 VGND VGND VPWR VPWR U$$184/A sky130_fd_sc_hd__a22o_1
XU$$194 U$$194/A U$$218/B VGND VGND VPWR VPWR U$$194/X sky130_fd_sc_hd__xor2_1
XFILLER_75_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_439 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_91_2 U$$3913/X U$$4046/X U$$4179/X VGND VGND VPWR VPWR dadda_fa_3_92_1/A
+ dadda_fa_3_91_3/A sky130_fd_sc_hd__fa_1
XFILLER_133_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1050 input82/X VGND VGND VPWR VPWR U$$3618/B1 sky130_fd_sc_hd__buf_6
Xrepeater1061 input81/X VGND VGND VPWR VPWR U$$3481/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_84_1 U$$4431/X input239/X dadda_fa_2_84_1/CIN VGND VGND VPWR VPWR dadda_fa_3_85_0/CIN
+ dadda_fa_3_84_2/CIN sky130_fd_sc_hd__fa_1
Xoutput258 output258/A VGND VGND VPWR VPWR o[100] sky130_fd_sc_hd__buf_2
XFILLER_173_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1072 input80/X VGND VGND VPWR VPWR U$$4027/A1 sky130_fd_sc_hd__buf_8
Xrepeater1083 U$$50/A1 VGND VGND VPWR VPWR U$$3749/A1 sky130_fd_sc_hd__buf_6
Xoutput269 output269/A VGND VGND VPWR VPWR o[110] sky130_fd_sc_hd__buf_2
Xdadda_fa_5_61_0 dadda_fa_5_61_0/A dadda_fa_5_61_0/B dadda_fa_5_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_62_0/A dadda_fa_6_61_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1094 U$$3882/B1 VGND VGND VPWR VPWR U$$48/A1 sky130_fd_sc_hd__buf_4
XFILLER_87_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_77_0 dadda_fa_2_77_0/A dadda_fa_2_77_0/B dadda_fa_2_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_0/B dadda_fa_3_77_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_60_8 dadda_fa_1_60_8/A dadda_fa_1_60_8/B dadda_fa_1_60_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_61_3/A dadda_fa_3_60_0/A sky130_fd_sc_hd__fa_2
XFILLER_67_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_53_7 U$$3172/X U$$3305/X U$$3438/X VGND VGND VPWR VPWR dadda_fa_2_54_2/CIN
+ dadda_fa_2_53_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_56_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1072 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_99_1 dadda_fa_4_99_1/A dadda_fa_4_99_1/B dadda_fa_4_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/B dadda_fa_5_99_1/B sky130_fd_sc_hd__fa_1
XFILLER_125_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_775 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_76_0 dadda_fa_7_76_0/A dadda_fa_7_76_0/B dadda_fa_7_76_0/CIN VGND VGND
+ VPWR VPWR _373_/D _244_/D sky130_fd_sc_hd__fa_1
XFILLER_180_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_948 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1043 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3208 U$$3208/A U$$3208/B VGND VGND VPWR VPWR U$$3208/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3219 U$$4452/A1 U$$3255/A2 U$$4454/A1 U$$3255/B2 VGND VGND VPWR VPWR U$$3220/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_282 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2507 U$$2507/A U$$2597/B VGND VGND VPWR VPWR U$$2507/X sky130_fd_sc_hd__xor2_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2518 U$$3612/B1 U$$2542/A2 U$$874/B1 U$$2542/B2 VGND VGND VPWR VPWR U$$2519/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2529 U$$2529/A U$$2577/B VGND VGND VPWR VPWR U$$2529/X sky130_fd_sc_hd__xor2_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1806 U$$1806/A U$$1840/B VGND VGND VPWR VPWR U$$1806/X sky130_fd_sc_hd__xor2_1
XU$$1817 U$$993/B1 U$$1819/A2 U$$860/A1 U$$1819/B2 VGND VGND VPWR VPWR U$$1818/A sky130_fd_sc_hd__a22o_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1828 U$$1828/A U$$1878/B VGND VGND VPWR VPWR U$$1828/X sky130_fd_sc_hd__xor2_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1839 U$$3618/B1 U$$1839/A2 U$$2113/B1 U$$1839/B2 VGND VGND VPWR VPWR U$$1840/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_324_ _325_/CLK _324_/D VGND VGND VPWR VPWR _324_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_255_ _255_/CLK _255_/D VGND VGND VPWR VPWR _255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_186_ _327_/CLK _186_/D VGND VGND VPWR VPWR _186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_94_0 dadda_fa_3_94_0/A dadda_fa_3_94_0/B dadda_fa_3_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_0/B dadda_fa_4_94_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater706 U$$3926/B2 VGND VGND VPWR VPWR U$$3946/B2 sky130_fd_sc_hd__buf_6
XFILLER_133_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater717 U$$3704/X VGND VGND VPWR VPWR U$$3777/B2 sky130_fd_sc_hd__buf_6
Xrepeater728 U$$3430/X VGND VGND VPWR VPWR U$$3479/B2 sky130_fd_sc_hd__buf_6
XFILLER_81_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4410 input128/X U$$4388/X U$$4410/B1 U$$4430/B2 VGND VGND VPWR VPWR U$$4411/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_56_5 dadda_fa_2_56_5/A dadda_fa_2_56_5/B dadda_fa_2_56_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_57_2/A dadda_fa_4_56_0/A sky130_fd_sc_hd__fa_1
XU$$4421 U$$4421/A U$$4421/B VGND VGND VPWR VPWR U$$4421/X sky130_fd_sc_hd__xor2_1
Xrepeater739 U$$3378/B2 VGND VGND VPWR VPWR U$$3390/B2 sky130_fd_sc_hd__buf_4
XU$$4432 U$$4432/A1 U$$4388/X U$$4434/A1 U$$4432/B2 VGND VGND VPWR VPWR U$$4433/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4431_1792 VGND VGND VPWR VPWR U$$4431_1792/HI U$$4431/B sky130_fd_sc_hd__conb_1
XU$$4443 U$$4443/A U$$4443/B VGND VGND VPWR VPWR U$$4443/X sky130_fd_sc_hd__xor2_1
XFILLER_64_111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4454 U$$4454/A1 U$$4388/X U$$4456/A1 U$$4498/B2 VGND VGND VPWR VPWR U$$4455/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_49_4 dadda_fa_2_49_4/A dadda_fa_2_49_4/B dadda_fa_2_49_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_1/CIN dadda_fa_3_49_3/CIN sky130_fd_sc_hd__fa_1
XU$$4465 U$$4465/A U$$4465/B VGND VGND VPWR VPWR U$$4465/X sky130_fd_sc_hd__xor2_1
XU$$3720 U$$3720/A U$$3740/B VGND VGND VPWR VPWR U$$3720/X sky130_fd_sc_hd__xor2_1
XU$$4476 U$$4476/A1 U$$4388/X U$$4476/B1 U$$4476/B2 VGND VGND VPWR VPWR U$$4477/A
+ sky130_fd_sc_hd__a22o_1
XU$$3731 U$$4277/B1 U$$3739/A2 U$$4418/A1 U$$3739/B2 VGND VGND VPWR VPWR U$$3732/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4487 U$$4487/A U$$4487/B VGND VGND VPWR VPWR U$$4487/X sky130_fd_sc_hd__xor2_1
XTAP_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3742 U$$3742/A U$$3778/B VGND VGND VPWR VPWR U$$3742/X sky130_fd_sc_hd__xor2_1
XTAP_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3753 input80/X U$$3753/A2 U$$4029/A1 U$$3753/B2 VGND VGND VPWR VPWR U$$3754/A
+ sky130_fd_sc_hd__a22o_1
XU$$4498 U$$4498/A1 U$$4388/X U$$4500/A1 U$$4498/B2 VGND VGND VPWR VPWR U$$4499/A
+ sky130_fd_sc_hd__a22o_1
XU$$3764 U$$3764/A U$$3774/B VGND VGND VPWR VPWR U$$3764/X sky130_fd_sc_hd__xor2_1
XFILLER_46_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3775 U$$3775/A1 U$$3703/X U$$3775/B1 U$$3704/X VGND VGND VPWR VPWR U$$3776/A sky130_fd_sc_hd__a22o_1
XU$$3786 U$$3786/A U$$3814/B VGND VGND VPWR VPWR U$$3786/X sky130_fd_sc_hd__xor2_1
XU$$4507_1830 VGND VGND VPWR VPWR U$$4507_1830/HI U$$4507/B sky130_fd_sc_hd__conb_1
XU$$3797 U$$4343/B1 U$$3813/A2 U$$4210/A1 U$$3813/B2 VGND VGND VPWR VPWR U$$3798/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_923 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_948 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_45_5 U$$2092/X U$$2225/X VGND VGND VPWR VPWR dadda_fa_2_46_3/CIN dadda_fa_3_45_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_87_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_51_4 U$$1705/X U$$1838/X U$$1971/X VGND VGND VPWR VPWR dadda_fa_2_52_1/CIN
+ dadda_fa_2_51_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$908 U$$84/B1 U$$918/A2 U$$910/A1 U$$918/B2 VGND VGND VPWR VPWR U$$909/A sky130_fd_sc_hd__a22o_1
XU$$919 U$$919/A U$$919/B VGND VGND VPWR VPWR U$$919/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_44_3 U$$1292/X U$$1425/X U$$1558/X VGND VGND VPWR VPWR dadda_fa_2_45_3/B
+ dadda_fa_2_44_5/B sky130_fd_sc_hd__fa_1
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_21_2 dadda_fa_4_21_2/A dadda_fa_4_21_2/B dadda_ha_3_21_3/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_22_0/CIN dadda_fa_5_21_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_14_1 U$$700/X U$$833/X U$$966/X VGND VGND VPWR VPWR dadda_fa_5_15_0/B
+ dadda_fa_5_14_1/B sky130_fd_sc_hd__fa_1
XFILLER_110_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_59_3 dadda_fa_3_59_3/A dadda_fa_3_59_3/B dadda_fa_3_59_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_60_1/B dadda_fa_4_59_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3005 U$$3416/A1 U$$3011/A2 input122/X U$$3011/B2 VGND VGND VPWR VPWR U$$3006/A
+ sky130_fd_sc_hd__a22o_1
XU$$3016 input40/X VGND VGND VPWR VPWR U$$3016/Y sky130_fd_sc_hd__inv_1
XU$$3027 U$$3027/A U$$3075/B VGND VGND VPWR VPWR U$$3027/X sky130_fd_sc_hd__xor2_1
XFILLER_189_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3038 input127/X U$$3124/A2 U$$26/A1 U$$3124/B2 VGND VGND VPWR VPWR U$$3039/A sky130_fd_sc_hd__a22o_1
XFILLER_90_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2304 U$$934/A1 U$$2308/A2 U$$936/A1 U$$2308/B2 VGND VGND VPWR VPWR U$$2305/A sky130_fd_sc_hd__a22o_1
XU$$3049 U$$3049/A U$$3083/B VGND VGND VPWR VPWR U$$3049/X sky130_fd_sc_hd__xor2_1
XU$$2315 U$$2315/A U$$2317/B VGND VGND VPWR VPWR U$$2315/X sky130_fd_sc_hd__xor2_1
XU$$2326 U$$956/A1 U$$2326/A2 U$$2326/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2327/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2337 U$$2609/B1 U$$2417/A2 U$$3296/B1 U$$2417/B2 VGND VGND VPWR VPWR U$$2338/A
+ sky130_fd_sc_hd__a22o_1
XU$$1603 U$$3108/B1 U$$1607/A2 U$$2975/A1 U$$1607/B2 VGND VGND VPWR VPWR U$$1604/A
+ sky130_fd_sc_hd__a22o_1
XU$$2348 U$$2348/A U$$2360/B VGND VGND VPWR VPWR U$$2348/X sky130_fd_sc_hd__xor2_1
XU$$1614 U$$1614/A U$$1628/B VGND VGND VPWR VPWR U$$1614/X sky130_fd_sc_hd__xor2_1
XFILLER_188_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2359 U$$3727/B1 U$$2359/A2 U$$4005/A1 U$$2359/B2 VGND VGND VPWR VPWR U$$2360/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_131_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1625 U$$4502/A1 U$$1637/A2 U$$2449/A1 U$$1637/B2 VGND VGND VPWR VPWR U$$1626/A
+ sky130_fd_sc_hd__a22o_1
XU$$1636 U$$1636/A U$$1638/B VGND VGND VPWR VPWR U$$1636/X sky130_fd_sc_hd__xor2_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1647 U$$1779/B U$$1647/B VGND VGND VPWR VPWR U$$1647/X sky130_fd_sc_hd__and2_1
XFILLER_61_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1658 U$$2343/A1 U$$1688/A2 U$$1932/B1 U$$1688/B2 VGND VGND VPWR VPWR U$$1659/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1669 U$$1669/A U$$1707/B VGND VGND VPWR VPWR U$$1669/X sky130_fd_sc_hd__xor2_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_307_ _327_/CLK _307_/D VGND VGND VPWR VPWR _307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_238_ _368_/CLK _238_/D VGND VGND VPWR VPWR _238_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_169_ _323_/CLK _169_/D VGND VGND VPWR VPWR _169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_61_3 dadda_fa_2_61_3/A dadda_fa_2_61_3/B dadda_fa_2_61_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/B dadda_fa_3_61_3/B sky130_fd_sc_hd__fa_1
Xrepeater503 U$$3098/A2 VGND VGND VPWR VPWR U$$3060/A2 sky130_fd_sc_hd__buf_4
XFILLER_38_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater514 U$$2949/A2 VGND VGND VPWR VPWR U$$2919/A2 sky130_fd_sc_hd__buf_6
XFILLER_97_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_2_108_0_1873 VGND VGND VPWR VPWR dadda_ha_2_108_0/A dadda_ha_2_108_0_1873/LO
+ sky130_fd_sc_hd__conb_1
Xrepeater525 U$$278/X VGND VGND VPWR VPWR U$$394/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_54_2 dadda_fa_2_54_2/A dadda_fa_2_54_2/B dadda_fa_2_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/A dadda_fa_3_54_3/A sky130_fd_sc_hd__fa_1
Xrepeater536 U$$2683/A2 VGND VGND VPWR VPWR U$$2625/A2 sky130_fd_sc_hd__clkbuf_4
Xrepeater547 U$$2524/A2 VGND VGND VPWR VPWR U$$2490/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater558 U$$2333/X VGND VGND VPWR VPWR U$$2449/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_5_31_1 dadda_fa_5_31_1/A dadda_fa_5_31_1/B dadda_fa_5_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_32_0/B dadda_fa_7_31_0/A sky130_fd_sc_hd__fa_1
XU$$4240 U$$4240/A1 U$$4240/A2 U$$4379/A1 U$$4240/B2 VGND VGND VPWR VPWR U$$4241/A
+ sky130_fd_sc_hd__a22o_1
XU$$4251 U$$4249/Y input59/X U$$4247/A U$$4250/X U$$4247/Y VGND VGND VPWR VPWR U$$4251/X
+ sky130_fd_sc_hd__a32o_4
Xrepeater569 U$$2099/A2 VGND VGND VPWR VPWR U$$2113/A2 sky130_fd_sc_hd__buf_4
XFILLER_26_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4262 U$$4262/A U$$4384/A VGND VGND VPWR VPWR U$$4262/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_47_1 U$$3160/X input198/X dadda_fa_2_47_1/CIN VGND VGND VPWR VPWR dadda_fa_3_48_0/CIN
+ dadda_fa_3_47_2/CIN sky130_fd_sc_hd__fa_1
XU$$4273 U$$4273/A1 U$$4275/A2 U$$4273/B1 U$$4275/B2 VGND VGND VPWR VPWR U$$4274/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4284 U$$4284/A U$$4370/B VGND VGND VPWR VPWR U$$4284/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_24_0 dadda_fa_5_24_0/A dadda_fa_5_24_0/B dadda_fa_5_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_25_0/A dadda_fa_6_24_0/CIN sky130_fd_sc_hd__fa_1
XU$$3550 U$$3550/A U$$3550/B VGND VGND VPWR VPWR U$$3550/X sky130_fd_sc_hd__xor2_1
XU$$4295 U$$4432/A1 U$$4297/A2 input78/X U$$4297/B2 VGND VGND VPWR VPWR U$$4296/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3561 U$$3561/A VGND VGND VPWR VPWR U$$3561/Y sky130_fd_sc_hd__inv_1
XU$$3572 U$$832/A1 U$$3660/A2 U$$3846/B1 U$$3660/B2 VGND VGND VPWR VPWR U$$3573/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3583 U$$3583/A U$$3609/B VGND VGND VPWR VPWR U$$3583/X sky130_fd_sc_hd__xor2_1
XU$$3594 U$$3594/A1 U$$3606/A2 U$$4005/B1 U$$3606/B2 VGND VGND VPWR VPWR U$$3595/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2860 U$$118/B1 U$$2868/A2 U$$122/A1 U$$2868/B2 VGND VGND VPWR VPWR U$$2861/A sky130_fd_sc_hd__a22o_1
XFILLER_34_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2871 U$$2871/A U$$2876/A VGND VGND VPWR VPWR U$$2871/X sky130_fd_sc_hd__xor2_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2882 U$$2880/B input36/X input37/X U$$2877/Y VGND VGND VPWR VPWR U$$2882/X sky130_fd_sc_hd__a22o_2
XU$$2893 U$$3987/B1 U$$2921/A2 U$$3852/B1 U$$2921/B2 VGND VGND VPWR VPWR U$$2894/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_1039 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1050 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1056 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_917 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_69_2 dadda_fa_4_69_2/A dadda_fa_4_69_2/B dadda_fa_4_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_70_0/CIN dadda_fa_5_69_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$800 final_adder.U$$800/A final_adder.U$$800/B VGND VGND VPWR VPWR
+ final_adder.U$$800/X sky130_fd_sc_hd__and2_1
XTAP_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_1_36_1 U$$478/X U$$611/X VGND VGND VPWR VPWR dadda_fa_2_37_5/B dadda_fa_3_36_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_102_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$811 final_adder.U$$778/A final_adder.U$$731/X final_adder.U$$699/X
+ VGND VGND VPWR VPWR final_adder.U$$811/X sky130_fd_sc_hd__a21o_1
XTAP_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_39_0 dadda_fa_7_39_0/A dadda_fa_7_39_0/B dadda_fa_7_39_0/CIN VGND VGND
+ VPWR VPWR _336_/D _207_/D sky130_fd_sc_hd__fa_2
XFILLER_112_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$833 final_adder.U$$800/A final_adder.U$$255/X final_adder.U$$721/X
+ VGND VGND VPWR VPWR final_adder.U$$833/X sky130_fd_sc_hd__a21o_1
XFILLER_25_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$855 final_adder.U$$758/X final_adder.U$$823/X final_adder.U$$759/X
+ VGND VGND VPWR VPWR final_adder.U$$855/X sky130_fd_sc_hd__a21o_2
XFILLER_186_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$705 U$$20/A1 U$$711/A2 U$$22/A1 U$$711/B2 VGND VGND VPWR VPWR U$$706/A sky130_fd_sc_hd__a22o_1
XFILLER_56_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$877 final_adder.U$$780/X final_adder.U$$733/X final_adder.U$$781/X
+ VGND VGND VPWR VPWR final_adder.U$$877/X sky130_fd_sc_hd__a21o_1
XFILLER_21_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$716 U$$716/A U$$740/B VGND VGND VPWR VPWR U$$716/X sky130_fd_sc_hd__xor2_1
XU$$727 U$$727/A1 U$$759/A2 U$$727/B1 U$$759/B2 VGND VGND VPWR VPWR U$$728/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_42_0 U$$91/X U$$224/X U$$357/X VGND VGND VPWR VPWR dadda_fa_2_43_3/A dadda_fa_2_42_4/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$738 U$$738/A U$$770/B VGND VGND VPWR VPWR U$$738/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$899 final_adder.U$$899/A1 final_adder.U$$837/X final_adder.U$$899/B1
+ VGND VGND VPWR VPWR final_adder.U$$899/X sky130_fd_sc_hd__a21o_1
XU$$749 U$$64/A1 U$$749/A2 U$$66/A1 U$$749/B2 VGND VGND VPWR VPWR U$$750/A sky130_fd_sc_hd__a22o_1
XFILLER_204_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_583 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1605 U$$930/B1 VGND VGND VPWR VPWR U$$932/A1 sky130_fd_sc_hd__buf_6
XFILLER_126_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1616 U$$4492/A1 VGND VGND VPWR VPWR U$$517/B1 sky130_fd_sc_hd__buf_6
XFILLER_192_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1627 input11/X VGND VGND VPWR VPWR U$$1370/A sky130_fd_sc_hd__buf_6
Xrepeater1638 input108/X VGND VGND VPWR VPWR U$$4077/B1 sky130_fd_sc_hd__buf_4
Xrepeater1649 U$$3116/B1 VGND VGND VPWR VPWR U$$2568/B1 sky130_fd_sc_hd__buf_6
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_71_2 dadda_fa_3_71_2/A dadda_fa_3_71_2/B dadda_fa_3_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_1/A dadda_fa_4_71_2/B sky130_fd_sc_hd__fa_1
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_64_1 dadda_fa_3_64_1/A dadda_fa_3_64_1/B dadda_fa_3_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_0/CIN dadda_fa_4_64_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_41_0 dadda_fa_6_41_0/A dadda_fa_6_41_0/B dadda_fa_6_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_42_0/B dadda_fa_7_41_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_57_0 dadda_fa_3_57_0/A dadda_fa_3_57_0/B dadda_fa_3_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_0/B dadda_fa_4_57_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2101 U$$44/B1 U$$2113/A2 U$$48/A1 U$$2113/B2 VGND VGND VPWR VPWR U$$2102/A sky130_fd_sc_hd__a22o_1
XU$$2112 U$$2112/A U$$2114/B VGND VGND VPWR VPWR U$$2112/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_100_2 dadda_fa_4_100_2/A dadda_fa_4_100_2/B dadda_fa_4_100_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_101_0/CIN dadda_fa_5_100_1/CIN sky130_fd_sc_hd__fa_1
XU$$2123 U$$2123/A1 U$$2149/A2 U$$616/B1 U$$2149/B2 VGND VGND VPWR VPWR U$$2124/A
+ sky130_fd_sc_hd__a22o_1
XU$$2134 U$$2134/A U$$2178/B VGND VGND VPWR VPWR U$$2134/X sky130_fd_sc_hd__xor2_1
XFILLER_62_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2145 U$$3102/B1 U$$2183/A2 U$$2967/B1 U$$2183/B2 VGND VGND VPWR VPWR U$$2146/A
+ sky130_fd_sc_hd__a22o_1
XU$$1400 U$$987/B1 U$$1404/A2 U$$854/A1 U$$1404/B2 VGND VGND VPWR VPWR U$$1401/A sky130_fd_sc_hd__a22o_1
XU$$1411 U$$1411/A U$$1423/B VGND VGND VPWR VPWR U$$1411/X sky130_fd_sc_hd__xor2_1
XU$$2156 U$$2156/A U$$2191/A VGND VGND VPWR VPWR U$$2156/X sky130_fd_sc_hd__xor2_1
XU$$1422 U$$461/B1 U$$1422/A2 U$$328/A1 U$$1422/B2 VGND VGND VPWR VPWR U$$1423/A sky130_fd_sc_hd__a22o_1
XFILLER_37_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2167 U$$934/A1 U$$2183/A2 U$$936/A1 U$$2183/B2 VGND VGND VPWR VPWR U$$2168/A sky130_fd_sc_hd__a22o_1
XFILLER_22_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1433 U$$1433/A U$$1459/B VGND VGND VPWR VPWR U$$1433/X sky130_fd_sc_hd__xor2_1
XU$$2178 U$$2178/A U$$2178/B VGND VGND VPWR VPWR U$$2178/X sky130_fd_sc_hd__xor2_1
XU$$2189 U$$3283/B1 U$$2189/A2 U$$2189/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2190/A
+ sky130_fd_sc_hd__a22o_1
XU$$1444 U$$2951/A1 U$$1448/A2 U$$1446/A1 U$$1448/B2 VGND VGND VPWR VPWR U$$1445/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1455 U$$1455/A U$$1501/B VGND VGND VPWR VPWR U$$1455/X sky130_fd_sc_hd__xor2_1
XU$$1466 U$$3108/B1 U$$1374/X U$$2975/A1 U$$1375/X VGND VGND VPWR VPWR U$$1467/A sky130_fd_sc_hd__a22o_1
XFILLER_203_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1477 U$$1477/A U$$1507/A VGND VGND VPWR VPWR U$$1477/X sky130_fd_sc_hd__xor2_1
XFILLER_188_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1488 U$$3680/A1 U$$1502/A2 U$$118/B1 U$$1502/B2 VGND VGND VPWR VPWR U$$1489/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1499 U$$1499/A U$$1499/B VGND VGND VPWR VPWR U$$1499/X sky130_fd_sc_hd__xor2_1
XFILLER_176_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_114_0 dadda_fa_7_114_0/A dadda_fa_7_114_0/B dadda_fa_7_114_0/CIN VGND
+ VGND VPWR VPWR _411_/D _282_/D sky130_fd_sc_hd__fa_1
XFILLER_30_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_79_1 dadda_fa_5_79_1/A dadda_fa_5_79_1/B dadda_fa_5_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_80_0/B dadda_fa_7_79_0/A sky130_fd_sc_hd__fa_1
XFILLER_143_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_951 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$107 _403_/Q _275_/Q VGND VGND VPWR VPWR final_adder.U$$149/B1 final_adder.U$$148/B
+ sky130_fd_sc_hd__ha_1
XFILLER_140_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$118 _414_/Q _286_/Q VGND VGND VPWR VPWR final_adder.U$$907/B1 final_adder.U$$136/A
+ sky130_fd_sc_hd__ha_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4070 U$$4070/A U$$4080/B VGND VGND VPWR VPWR U$$4070/X sky130_fd_sc_hd__xor2_1
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater388 U$$1057/A2 VGND VGND VPWR VPWR U$$997/A2 sky130_fd_sc_hd__buf_4
XU$$4081 U$$517/B1 U$$4103/A2 U$$384/A1 U$$4103/B2 VGND VGND VPWR VPWR U$$4082/A sky130_fd_sc_hd__a22o_1
Xrepeater399 U$$826/X VGND VGND VPWR VPWR U$$938/A2 sky130_fd_sc_hd__buf_4
XFILLER_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4092 U$$4092/A U$$4110/A VGND VGND VPWR VPWR U$$4092/X sky130_fd_sc_hd__xor2_1
XFILLER_25_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3380 U$$3517/A1 U$$3388/A2 input102/X U$$3390/B2 VGND VGND VPWR VPWR U$$3381/A
+ sky130_fd_sc_hd__a22o_1
XU$$3391 U$$3391/A U$$3395/B VGND VGND VPWR VPWR U$$3391/X sky130_fd_sc_hd__xor2_1
XFILLER_81_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2690 U$$2690/A U$$2739/A VGND VGND VPWR VPWR U$$2690/X sky130_fd_sc_hd__xor2_1
XFILLER_34_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_81_1 dadda_fa_4_81_1/A dadda_fa_4_81_1/B dadda_fa_4_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/B dadda_fa_5_81_1/B sky130_fd_sc_hd__fa_1
XFILLER_135_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_74_0 dadda_fa_4_74_0/A dadda_fa_4_74_0/B dadda_fa_4_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/A dadda_fa_5_74_1/A sky130_fd_sc_hd__fa_1
XFILLER_89_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput103 b[44] VGND VGND VPWR VPWR input103/X sky130_fd_sc_hd__buf_6
XFILLER_163_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput114 b[54] VGND VGND VPWR VPWR input114/X sky130_fd_sc_hd__buf_6
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput125 b[6] VGND VGND VPWR VPWR input125/X sky130_fd_sc_hd__buf_6
XTAP_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput136 c[106] VGND VGND VPWR VPWR input136/X sky130_fd_sc_hd__buf_4
XTAP_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput147 c[116] VGND VGND VPWR VPWR input147/X sky130_fd_sc_hd__clkbuf_4
XTAP_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput158 c[126] VGND VGND VPWR VPWR input158/X sky130_fd_sc_hd__clkbuf_2
XTAP_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput169 c[20] VGND VGND VPWR VPWR input169/X sky130_fd_sc_hd__clkbuf_4
Xfinal_adder.U$$630 final_adder.U$$646/B final_adder.U$$630/B VGND VGND VPWR VPWR
+ final_adder.U$$742/B sky130_fd_sc_hd__and2_1
XTAP_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$641 final_adder.U$$640/B final_adder.U$$537/X final_adder.U$$521/X
+ VGND VGND VPWR VPWR final_adder.U$$641/X sky130_fd_sc_hd__a21o_1
XTAP_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$652 final_adder.U$$668/B final_adder.U$$652/B VGND VGND VPWR VPWR
+ final_adder.U$$764/B sky130_fd_sc_hd__and2_1
XTAP_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$663 final_adder.U$$662/B final_adder.U$$559/X final_adder.U$$543/X
+ VGND VGND VPWR VPWR final_adder.U$$663/X sky130_fd_sc_hd__a21o_1
XTAP_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$502 U$$502/A U$$504/B VGND VGND VPWR VPWR U$$502/X sky130_fd_sc_hd__xor2_1
XFILLER_91_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$674 final_adder.U$$690/B final_adder.U$$674/B VGND VGND VPWR VPWR
+ final_adder.U$$786/B sky130_fd_sc_hd__and2_1
XU$$513 U$$650/A1 U$$515/A2 U$$652/A1 U$$515/B2 VGND VGND VPWR VPWR U$$514/A sky130_fd_sc_hd__a22o_1
XTAP_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$685 final_adder.U$$684/B final_adder.U$$581/X final_adder.U$$565/X
+ VGND VGND VPWR VPWR final_adder.U$$685/X sky130_fd_sc_hd__a21o_1
XTAP_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$524 U$$524/A U$$546/B VGND VGND VPWR VPWR U$$524/X sky130_fd_sc_hd__xor2_1
XFILLER_205_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$696 final_adder.U$$712/B final_adder.U$$696/B VGND VGND VPWR VPWR
+ final_adder.U$$776/A sky130_fd_sc_hd__and2_1
XTAP_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$535 U$$807/B1 U$$537/A2 U$$674/A1 U$$537/B2 VGND VGND VPWR VPWR U$$536/A sky130_fd_sc_hd__a22o_1
XFILLER_205_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$546 U$$546/A U$$546/B VGND VGND VPWR VPWR U$$546/X sky130_fd_sc_hd__xor2_1
XFILLER_189_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$557 U$$557/A U$$579/B VGND VGND VPWR VPWR U$$557/X sky130_fd_sc_hd__xor2_1
XTAP_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$568 U$$20/A1 U$$578/A2 U$$842/B1 U$$578/B2 VGND VGND VPWR VPWR U$$569/A sky130_fd_sc_hd__a22o_1
XU$$579 U$$579/A U$$579/B VGND VGND VPWR VPWR U$$579/X sky130_fd_sc_hd__xor2_1
XFILLER_112_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_386 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_89_0 dadda_fa_6_89_0/A dadda_fa_6_89_0/B dadda_fa_6_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_90_0/B dadda_fa_7_89_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1402 U$$2184/B VGND VGND VPWR VPWR U$$2191/A sky130_fd_sc_hd__buf_6
Xrepeater1413 U$$1991/B VGND VGND VPWR VPWR U$$1971/B sky130_fd_sc_hd__buf_8
XFILLER_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1424 U$$1914/B VGND VGND VPWR VPWR U$$1880/B sky130_fd_sc_hd__buf_6
Xrepeater1435 U$$1780/A VGND VGND VPWR VPWR U$$1751/B sky130_fd_sc_hd__buf_8
Xrepeater1446 input16/X VGND VGND VPWR VPWR U$$1644/A sky130_fd_sc_hd__buf_4
XFILLER_181_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1457 U$$983/B1 VGND VGND VPWR VPWR U$$846/B1 sky130_fd_sc_hd__buf_4
Xrepeater1468 U$$3584/B1 VGND VGND VPWR VPWR U$$709/A1 sky130_fd_sc_hd__buf_6
XFILLER_207_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1479 input126/X VGND VGND VPWR VPWR U$$842/B1 sky130_fd_sc_hd__buf_4
XFILLER_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1230 U$$1504/A1 U$$1230/A2 U$$1230/B1 U$$1230/B2 VGND VGND VPWR VPWR U$$1231/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1241 U$$1515/A1 U$$1311/A2 U$$969/A1 U$$1271/B2 VGND VGND VPWR VPWR U$$1242/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1252 U$$1252/A U$$1270/B VGND VGND VPWR VPWR U$$1252/X sky130_fd_sc_hd__xor2_1
XU$$1263 U$$987/B1 U$$1271/A2 U$$854/A1 U$$1281/B2 VGND VGND VPWR VPWR U$$1264/A sky130_fd_sc_hd__a22o_1
XFILLER_176_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1274 U$$1274/A U$$1316/B VGND VGND VPWR VPWR U$$1274/X sky130_fd_sc_hd__xor2_1
XU$$1285 U$$461/B1 U$$1289/A2 U$$328/A1 U$$1291/B2 VGND VGND VPWR VPWR U$$1286/A sky130_fd_sc_hd__a22o_1
XFILLER_203_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1296 U$$1296/A U$$1354/B VGND VGND VPWR VPWR U$$1296/X sky130_fd_sc_hd__xor2_1
XFILLER_31_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_91_0 dadda_fa_5_91_0/A dadda_fa_5_91_0/B dadda_fa_5_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_92_0/A dadda_fa_6_91_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_50_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1075 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1090 final_adder.U$$188/A final_adder.U$$897/X VGND VGND VPWR VPWR
+ output347/A sky130_fd_sc_hd__xor2_1
XFILLER_131_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_76_6 U$$3883/X U$$4016/X U$$4149/X VGND VGND VPWR VPWR dadda_fa_2_77_2/B
+ dadda_fa_2_76_5/B sky130_fd_sc_hd__fa_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_69_5 U$$4401/X input222/X dadda_fa_1_69_5/CIN VGND VGND VPWR VPWR dadda_fa_2_70_2/A
+ dadda_fa_2_69_5/A sky130_fd_sc_hd__fa_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _200_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_219 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_426 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_96_0 dadda_ha_1_96_0/A U$$2327/X VGND VGND VPWR VPWR dadda_fa_3_97_0/A
+ dadda_fa_3_96_0/A sky130_fd_sc_hd__ha_1
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_100_1 dadda_fa_3_100_1/A dadda_fa_3_100_1/B dadda_fa_3_100_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_0/CIN dadda_fa_4_100_2/A sky130_fd_sc_hd__fa_1
XFILLER_101_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_121_0 dadda_fa_6_121_0/A dadda_fa_6_121_0/B dadda_fa_6_121_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_122_0/B dadda_fa_7_121_0/CIN sky130_fd_sc_hd__fa_1
XTAP_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1099 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_64_4 U$$1731/X U$$1864/X U$$1997/X VGND VGND VPWR VPWR dadda_fa_1_65_6/CIN
+ dadda_fa_1_64_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_40_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_41_3 dadda_fa_3_41_3/A dadda_fa_3_41_3/B dadda_fa_3_41_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_42_1/B dadda_fa_4_41_2/CIN sky130_fd_sc_hd__fa_1
XTAP_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$460 final_adder.U$$464/B final_adder.U$$460/B VGND VGND VPWR VPWR
+ final_adder.U$$584/B sky130_fd_sc_hd__and2_1
XTAP_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$471 final_adder.U$$470/B final_adder.U$$349/X final_adder.U$$345/X
+ VGND VGND VPWR VPWR final_adder.U$$471/X sky130_fd_sc_hd__a21o_1
XTAP_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$310 U$$719/B1 U$$340/A2 U$$312/A1 U$$340/B2 VGND VGND VPWR VPWR U$$311/A sky130_fd_sc_hd__a22o_1
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$482 final_adder.U$$486/B final_adder.U$$482/B VGND VGND VPWR VPWR
+ final_adder.U$$606/B sky130_fd_sc_hd__and2_1
XTAP_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$321 U$$321/A U$$351/B VGND VGND VPWR VPWR U$$321/X sky130_fd_sc_hd__xor2_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_34_2 dadda_fa_3_34_2/A dadda_fa_3_34_2/B dadda_fa_3_34_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_1/A dadda_fa_4_34_2/B sky130_fd_sc_hd__fa_1
XTAP_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$493 final_adder.U$$492/B final_adder.U$$371/X final_adder.U$$367/X
+ VGND VGND VPWR VPWR final_adder.U$$493/X sky130_fd_sc_hd__a21o_1
XTAP_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$332 U$$56/B1 U$$350/A2 U$$882/A1 U$$350/B2 VGND VGND VPWR VPWR U$$333/A sky130_fd_sc_hd__a22o_1
XTAP_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$343 U$$343/A U$$343/B VGND VGND VPWR VPWR U$$343/X sky130_fd_sc_hd__xor2_1
XFILLER_189_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$354 U$$763/B1 U$$396/A2 U$$630/A1 U$$396/B2 VGND VGND VPWR VPWR U$$355/A sky130_fd_sc_hd__a22o_1
XTAP_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$365 U$$365/A U$$397/B VGND VGND VPWR VPWR U$$365/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_27_1 U$$1524/X U$$1657/X U$$1790/X VGND VGND VPWR VPWR dadda_fa_4_28_0/CIN
+ dadda_fa_4_27_2/A sky130_fd_sc_hd__fa_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$376 U$$650/A1 U$$378/A2 U$$652/A1 U$$378/B2 VGND VGND VPWR VPWR U$$377/A sky130_fd_sc_hd__a22o_1
XU$$387 U$$387/A U$$395/B VGND VGND VPWR VPWR U$$387/X sky130_fd_sc_hd__xor2_1
XU$$398 U$$807/B1 U$$278/X U$$674/A1 U$$279/X VGND VGND VPWR VPWR U$$399/A sky130_fd_sc_hd__a22o_1
XFILLER_177_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1004 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_954 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1210 U$$625/B VGND VGND VPWR VPWR U$$617/B sky130_fd_sc_hd__buf_6
Xrepeater1221 U$$546/B VGND VGND VPWR VPWR U$$528/B sky130_fd_sc_hd__buf_8
XFILLER_160_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1232 U$$4165/B VGND VGND VPWR VPWR U$$4145/B sky130_fd_sc_hd__buf_6
Xrepeater1243 U$$343/B VGND VGND VPWR VPWR U$$317/B sky130_fd_sc_hd__buf_4
XFILLER_181_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1254 U$$4044/B VGND VGND VPWR VPWR U$$4036/B sky130_fd_sc_hd__buf_8
Xdadda_fa_2_86_5 dadda_fa_2_86_5/A dadda_fa_2_86_5/B dadda_fa_2_86_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_87_2/A dadda_fa_4_86_0/A sky130_fd_sc_hd__fa_2
Xrepeater1265 U$$3971/B VGND VGND VPWR VPWR U$$3909/B sky130_fd_sc_hd__buf_8
XFILLER_126_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1276 U$$919/B VGND VGND VPWR VPWR U$$847/B sky130_fd_sc_hd__buf_6
Xrepeater1287 U$$3623/B VGND VGND VPWR VPWR U$$3665/B sky130_fd_sc_hd__buf_6
XFILLER_113_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1298 U$$3518/B VGND VGND VPWR VPWR U$$3490/B sky130_fd_sc_hd__buf_6
XFILLER_141_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_79_4 dadda_fa_2_79_4/A dadda_fa_2_79_4/B dadda_fa_2_79_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_1/CIN dadda_fa_3_79_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1060 U$$1060/A U$$1076/B VGND VGND VPWR VPWR U$$1060/X sky130_fd_sc_hd__xor2_1
XFILLER_195_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1071 U$$932/B1 U$$963/X U$$799/A1 U$$964/X VGND VGND VPWR VPWR U$$1072/A sky130_fd_sc_hd__a22o_1
XFILLER_51_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1082 U$$1082/A U$$1095/A VGND VGND VPWR VPWR U$$1082/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1093 U$$1504/A1 U$$1093/A2 U$$1093/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1094/A
+ sky130_fd_sc_hd__a22o_1
XU$$3157_1745 VGND VGND VPWR VPWR U$$3157_1745/HI U$$3157/A1 sky130_fd_sc_hd__conb_1
XFILLER_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_116_1 dadda_fa_5_116_1/A dadda_fa_5_116_1/B dadda_fa_5_116_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_117_0/B dadda_fa_7_116_0/A sky130_fd_sc_hd__fa_1
XFILLER_192_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_109_0 dadda_fa_5_109_0/A dadda_fa_5_109_0/B dadda_fa_5_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_110_0/A dadda_fa_6_109_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_81_4 U$$2829/X U$$2962/X U$$3095/X VGND VGND VPWR VPWR dadda_fa_2_82_2/B
+ dadda_fa_2_81_5/A sky130_fd_sc_hd__fa_1
XFILLER_63_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_74_3 U$$2948/X U$$3081/X U$$3214/X VGND VGND VPWR VPWR dadda_fa_2_75_1/B
+ dadda_fa_2_74_4/B sky130_fd_sc_hd__fa_1
XFILLER_98_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_51_2 dadda_fa_4_51_2/A dadda_fa_4_51_2/B dadda_fa_4_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_52_0/CIN dadda_fa_5_51_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_67_2 U$$3333/X U$$3466/X U$$3599/X VGND VGND VPWR VPWR dadda_fa_2_68_1/A
+ dadda_fa_2_67_4/A sky130_fd_sc_hd__fa_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_44_1 dadda_fa_4_44_1/A dadda_fa_4_44_1/B dadda_fa_4_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/B dadda_fa_5_44_1/B sky130_fd_sc_hd__fa_1
XFILLER_86_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_21_0 dadda_fa_7_21_0/A dadda_fa_7_21_0/B dadda_fa_7_21_0/CIN VGND VGND
+ VPWR VPWR _318_/D _189_/D sky130_fd_sc_hd__fa_1
XFILLER_73_315 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_37_0 dadda_fa_4_37_0/A dadda_fa_4_37_0/B dadda_fa_4_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/A dadda_fa_5_37_1/A sky130_fd_sc_hd__fa_1
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_340_ _342_/CLK _340_/D VGND VGND VPWR VPWR _340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_271_ _394_/CLK _271_/D VGND VGND VPWR VPWR _271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_751 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_70_4 U$$2009/X U$$2142/X VGND VGND VPWR VPWR dadda_fa_1_71_7/CIN dadda_fa_2_70_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_182_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_89_3 dadda_fa_3_89_3/A dadda_fa_3_89_3/B dadda_fa_3_89_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_90_1/B dadda_fa_4_89_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_0_56_2 U$$917/X U$$1050/X VGND VGND VPWR VPWR dadda_fa_1_57_8/A dadda_fa_2_56_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_111_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_62_1 U$$530/X U$$663/X U$$796/X VGND VGND VPWR VPWR dadda_fa_1_63_5/CIN
+ dadda_fa_1_62_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_209_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3902 U$$4176/A1 U$$3902/A2 U$$3902/B1 U$$3902/B2 VGND VGND VPWR VPWR U$$3903/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_55_0 U$$117/X U$$250/X U$$383/X VGND VGND VPWR VPWR dadda_fa_1_56_7/CIN
+ dadda_fa_1_55_8/CIN sky130_fd_sc_hd__fa_1
XU$$3913 U$$3913/A U$$3967/B VGND VGND VPWR VPWR U$$3913/X sky130_fd_sc_hd__xor2_1
XU$$3924 U$$4333/B1 U$$3926/A2 U$$912/A1 U$$3926/B2 VGND VGND VPWR VPWR U$$3925/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3935 U$$3935/A U$$3947/B VGND VGND VPWR VPWR U$$3935/X sky130_fd_sc_hd__xor2_1
XTAP_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3946 U$$384/A1 U$$3946/A2 U$$3946/B1 U$$3946/B2 VGND VGND VPWR VPWR U$$3947/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3957 U$$3957/A U$$3972/A VGND VGND VPWR VPWR U$$3957/X sky130_fd_sc_hd__xor2_1
XTAP_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$290 final_adder.U$$292/B final_adder.U$$290/B VGND VGND VPWR VPWR
+ final_adder.U$$416/B sky130_fd_sc_hd__and2_1
XTAP_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3968 U$$4379/A1 U$$3968/A2 input124/X U$$3968/B2 VGND VGND VPWR VPWR U$$3969/A
+ sky130_fd_sc_hd__a22o_1
XU$$140 U$$272/B U$$140/B VGND VGND VPWR VPWR U$$140/X sky130_fd_sc_hd__and2_1
XFILLER_91_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$151 U$$14/A1 U$$175/A2 U$$16/A1 U$$175/B2 VGND VGND VPWR VPWR U$$152/A sky130_fd_sc_hd__a22o_1
XFILLER_17_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3979 U$$3979/A1 U$$4011/A2 U$$3979/B1 U$$4011/B2 VGND VGND VPWR VPWR U$$3980/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$162 U$$162/A U$$184/B VGND VGND VPWR VPWR U$$162/X sky130_fd_sc_hd__xor2_1
XTAP_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$173 U$$36/A1 U$$175/A2 U$$38/A1 U$$175/B2 VGND VGND VPWR VPWR U$$174/A sky130_fd_sc_hd__a22o_1
XFILLER_150_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$184 U$$184/A U$$184/B VGND VGND VPWR VPWR U$$184/X sky130_fd_sc_hd__xor2_1
XU$$195 U$$58/A1 U$$217/A2 U$$60/A1 U$$217/B2 VGND VGND VPWR VPWR U$$196/A sky130_fd_sc_hd__a22o_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4425_1789 VGND VGND VPWR VPWR U$$4425_1789/HI U$$4425/B sky130_fd_sc_hd__conb_1
XFILLER_207_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_91_3 U$$4312/X U$$4445/X input247/X VGND VGND VPWR VPWR dadda_fa_3_92_1/B
+ dadda_fa_3_91_3/B sky130_fd_sc_hd__fa_1
XFILLER_114_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1040 U$$3483/B1 VGND VGND VPWR VPWR U$$745/A1 sky130_fd_sc_hd__buf_4
XFILLER_142_832 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1051 input82/X VGND VGND VPWR VPWR U$$741/B1 sky130_fd_sc_hd__buf_6
XFILLER_5_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_84_2 dadda_fa_2_84_2/A dadda_fa_2_84_2/B dadda_fa_2_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/A dadda_fa_3_84_3/A sky130_fd_sc_hd__fa_1
XU$$2061_1727 VGND VGND VPWR VPWR U$$2061_1727/HI U$$2061/A1 sky130_fd_sc_hd__conb_1
Xrepeater1062 input81/X VGND VGND VPWR VPWR U$$3344/A1 sky130_fd_sc_hd__buf_8
Xoutput259 output259/A VGND VGND VPWR VPWR o[101] sky130_fd_sc_hd__buf_2
Xrepeater1073 input79/X VGND VGND VPWR VPWR U$$3749/B1 sky130_fd_sc_hd__buf_6
Xrepeater1084 U$$2925/B1 VGND VGND VPWR VPWR U$$461/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_61_1 dadda_fa_5_61_1/A dadda_fa_5_61_1/B dadda_fa_5_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_62_0/B dadda_fa_7_61_0/A sky130_fd_sc_hd__fa_2
XFILLER_102_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1095 U$$3747/A1 VGND VGND VPWR VPWR U$$3882/B1 sky130_fd_sc_hd__buf_8
Xdadda_fa_2_77_1 dadda_fa_2_77_1/A dadda_fa_2_77_1/B dadda_fa_2_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_0/CIN dadda_fa_3_77_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_54_0 dadda_fa_5_54_0/A dadda_fa_5_54_0/B dadda_fa_5_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_55_0/A dadda_fa_6_54_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_136_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_53_8 U$$3571/X input205/X dadda_fa_1_53_8/CIN VGND VGND VPWR VPWR dadda_fa_2_54_3/A
+ dadda_fa_3_53_0/A sky130_fd_sc_hd__fa_1
XFILLER_82_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_100_0 dadda_fa_2_100_0/A U$$2601/X U$$2734/X VGND VGND VPWR VPWR dadda_fa_3_101_1/B
+ dadda_fa_3_100_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_51_532 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_99_2 dadda_fa_4_99_2/A dadda_fa_4_99_2/B dadda_fa_4_99_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_100_0/CIN dadda_fa_5_99_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_180_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_69_0 dadda_fa_7_69_0/A dadda_fa_7_69_0/B dadda_fa_7_69_0/CIN VGND VGND
+ VPWR VPWR _366_/D _237_/D sky130_fd_sc_hd__fa_1
XFILLER_105_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_72_0 U$$2013/X U$$2146/X U$$2279/X VGND VGND VPWR VPWR dadda_fa_2_73_0/B
+ dadda_fa_2_72_3/B sky130_fd_sc_hd__fa_1
XFILLER_28_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_1153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3209 U$$741/B1 U$$3229/A2 U$$3485/A1 U$$3227/B2 VGND VGND VPWR VPWR U$$3210/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2508 U$$4013/B1 U$$2596/A2 U$$4015/B1 U$$2596/B2 VGND VGND VPWR VPWR U$$2509/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2519 U$$2519/A U$$2543/B VGND VGND VPWR VPWR U$$2519/X sky130_fd_sc_hd__xor2_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1807 U$$2901/B1 U$$1831/A2 U$$4410/B1 U$$1831/B2 VGND VGND VPWR VPWR U$$1808/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1818 U$$1818/A U$$1820/B VGND VGND VPWR VPWR U$$1818/X sky130_fd_sc_hd__xor2_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_746 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1829 U$$594/B1 U$$1831/A2 U$$598/A1 U$$1831/B2 VGND VGND VPWR VPWR U$$1830/A sky130_fd_sc_hd__a22o_1
XFILLER_199_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_323_ _323_/CLK _323_/D VGND VGND VPWR VPWR _323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_254_ _382_/CLK _254_/D VGND VGND VPWR VPWR _254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_185_ _314_/CLK _185_/D VGND VGND VPWR VPWR _185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_94_1 dadda_fa_3_94_1/A dadda_fa_3_94_1/B dadda_fa_3_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_0/CIN dadda_fa_4_94_2/A sky130_fd_sc_hd__fa_1
XFILLER_182_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_71_0 dadda_fa_6_71_0/A dadda_fa_6_71_0/B dadda_fa_6_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_72_0/B dadda_fa_7_71_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_87_0 dadda_fa_3_87_0/A dadda_fa_3_87_0/B dadda_fa_3_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_0/B dadda_fa_4_87_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater707 U$$3966/B2 VGND VGND VPWR VPWR U$$3926/B2 sky130_fd_sc_hd__buf_6
XU$$4400 U$$4400/A1 U$$4388/X U$$4402/A1 U$$4432/B2 VGND VGND VPWR VPWR U$$4401/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater718 U$$3612/B2 VGND VGND VPWR VPWR U$$3606/B2 sky130_fd_sc_hd__buf_6
Xrepeater729 U$$3489/B2 VGND VGND VPWR VPWR U$$3527/B2 sky130_fd_sc_hd__buf_6
XFILLER_133_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4411 U$$4411/A U$$4411/B VGND VGND VPWR VPWR U$$4411/X sky130_fd_sc_hd__xor2_1
XU$$4422 U$$4422/A1 U$$4388/X U$$4424/A1 U$$4426/B2 VGND VGND VPWR VPWR U$$4423/A
+ sky130_fd_sc_hd__a22o_1
XU$$4433 U$$4433/A U$$4433/B VGND VGND VPWR VPWR U$$4433/X sky130_fd_sc_hd__xor2_1
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4444 input83/X U$$4388/X input84/X U$$4498/B2 VGND VGND VPWR VPWR U$$4445/A sky130_fd_sc_hd__a22o_1
XU$$3710 U$$3710/A U$$3794/B VGND VGND VPWR VPWR U$$3710/X sky130_fd_sc_hd__xor2_1
XU$$4455 U$$4455/A U$$4455/B VGND VGND VPWR VPWR U$$4455/X sky130_fd_sc_hd__xor2_1
XFILLER_92_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4466 U$$4466/A1 U$$4388/X U$$4466/B1 U$$4476/B2 VGND VGND VPWR VPWR U$$4467/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_116_0 U$$3830/X U$$3963/X U$$4096/X VGND VGND VPWR VPWR dadda_fa_5_117_0/A
+ dadda_fa_5_116_1/A sky130_fd_sc_hd__fa_1
XU$$3721 U$$4269/A1 U$$3739/A2 U$$4269/B1 U$$3739/B2 VGND VGND VPWR VPWR U$$3722/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_49_5 dadda_fa_2_49_5/A dadda_fa_2_49_5/B dadda_fa_2_49_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_50_2/A dadda_fa_4_49_0/A sky130_fd_sc_hd__fa_2
XTAP_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4477 U$$4477/A U$$4477/B VGND VGND VPWR VPWR U$$4477/X sky130_fd_sc_hd__xor2_1
XTAP_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3732 U$$3732/A U$$3740/B VGND VGND VPWR VPWR U$$3732/X sky130_fd_sc_hd__xor2_1
XU$$4488 U$$4488/A1 U$$4388/X U$$4490/A1 U$$4494/B2 VGND VGND VPWR VPWR U$$4489/A
+ sky130_fd_sc_hd__a22o_1
XU$$3743 U$$4428/A1 U$$3777/A2 input75/X U$$3777/B2 VGND VGND VPWR VPWR U$$3744/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4499 U$$4499/A U$$4499/B VGND VGND VPWR VPWR U$$4499/X sky130_fd_sc_hd__xor2_1
XU$$3754 U$$3754/A U$$3754/B VGND VGND VPWR VPWR U$$3754/X sky130_fd_sc_hd__xor2_1
XU$$3765 U$$4176/A1 U$$3773/A2 U$$3902/B1 U$$3773/B2 VGND VGND VPWR VPWR U$$3766/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3776 U$$3776/A U$$3836/A VGND VGND VPWR VPWR U$$3776/X sky130_fd_sc_hd__xor2_1
XTAP_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3787 U$$3922/B1 U$$3793/A2 U$$3787/B1 U$$3793/B2 VGND VGND VPWR VPWR U$$3788/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3798 U$$3798/A U$$3814/B VGND VGND VPWR VPWR U$$3798/X sky130_fd_sc_hd__xor2_1
XFILLER_61_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_692 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_28 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_51_5 U$$2104/X U$$2237/X U$$2370/X VGND VGND VPWR VPWR dadda_fa_2_52_2/A
+ dadda_fa_2_51_5/A sky130_fd_sc_hd__fa_1
XFILLER_96_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$909 U$$909/A U$$919/B VGND VGND VPWR VPWR U$$909/X sky130_fd_sc_hd__xor2_1
XFILLER_55_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_44_4 U$$1691/X U$$1824/X U$$1957/X VGND VGND VPWR VPWR dadda_fa_2_45_3/CIN
+ dadda_fa_2_44_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_37_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_14_2 U$$968/B input162/X dadda_ha_3_14_0/SUM VGND VGND VPWR VPWR dadda_fa_5_15_0/CIN
+ dadda_fa_5_14_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_145_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_104_0_1862 VGND VGND VPWR VPWR dadda_fa_2_104_0/A dadda_fa_2_104_0_1862/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_106_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_832 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3006 U$$3006/A U$$3013/A VGND VGND VPWR VPWR U$$3006/X sky130_fd_sc_hd__xor2_1
XFILLER_115_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3017 input40/X U$$3017/B VGND VGND VPWR VPWR U$$3017/X sky130_fd_sc_hd__and2_1
XU$$3028 U$$3028/A1 U$$3060/A2 U$$3987/B1 U$$3060/B2 VGND VGND VPWR VPWR U$$3029/A
+ sky130_fd_sc_hd__a22o_1
XU$$3039 U$$3039/A U$$3125/B VGND VGND VPWR VPWR U$$3039/X sky130_fd_sc_hd__xor2_1
XFILLER_207_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2305 U$$2305/A U$$2309/B VGND VGND VPWR VPWR U$$2305/X sky130_fd_sc_hd__xor2_1
XFILLER_46_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2316 U$$2316/A1 U$$2316/A2 U$$4236/A1 U$$2316/B2 VGND VGND VPWR VPWR U$$2317/A
+ sky130_fd_sc_hd__a22o_1
XU$$2327 U$$2327/A U$$2328/A VGND VGND VPWR VPWR U$$2327/X sky130_fd_sc_hd__xor2_1
XU$$2338 U$$2338/A U$$2366/B VGND VGND VPWR VPWR U$$2338/X sky130_fd_sc_hd__xor2_1
XU$$2349 U$$2623/A1 U$$2359/A2 U$$2625/A1 U$$2359/B2 VGND VGND VPWR VPWR U$$2350/A
+ sky130_fd_sc_hd__a22o_1
XU$$1604 U$$1604/A U$$1608/B VGND VGND VPWR VPWR U$$1604/X sky130_fd_sc_hd__xor2_1
XFILLER_76_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1615 U$$930/A1 U$$1635/A2 U$$2165/A1 U$$1635/B2 VGND VGND VPWR VPWR U$$1616/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1626 U$$1626/A U$$1638/B VGND VGND VPWR VPWR U$$1626/X sky130_fd_sc_hd__xor2_1
XFILLER_188_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1637 U$$4514/A1 U$$1637/A2 U$$4516/A1 U$$1637/B2 VGND VGND VPWR VPWR U$$1638/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1648 U$$1646/Y input17/X U$$1644/A U$$1647/X U$$1644/Y VGND VGND VPWR VPWR U$$1648/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_202_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1659 U$$1659/A U$$1689/B VGND VGND VPWR VPWR U$$1659/X sky130_fd_sc_hd__xor2_1
XFILLER_42_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_306_ _326_/CLK _306_/D VGND VGND VPWR VPWR _306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_721 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_237_ _367_/CLK _237_/D VGND VGND VPWR VPWR _237_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_168_ _325_/CLK _168_/D VGND VGND VPWR VPWR _168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_61_4 dadda_fa_2_61_4/A dadda_fa_2_61_4/B dadda_fa_2_61_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_1/CIN dadda_fa_3_61_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_85_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater504 U$$3098/A2 VGND VGND VPWR VPWR U$$3108/A2 sky130_fd_sc_hd__buf_6
XFILLER_85_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater515 U$$2967/A2 VGND VGND VPWR VPWR U$$2949/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater526 U$$278/X VGND VGND VPWR VPWR U$$396/A2 sky130_fd_sc_hd__buf_4
XFILLER_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_54_3 dadda_fa_2_54_3/A dadda_fa_2_54_3/B dadda_fa_2_54_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/B dadda_fa_3_54_3/B sky130_fd_sc_hd__fa_1
Xrepeater537 U$$2683/A2 VGND VGND VPWR VPWR U$$2653/A2 sky130_fd_sc_hd__buf_4
XU$$4230 U$$4504/A1 U$$4240/A2 U$$4506/A1 U$$4240/B2 VGND VGND VPWR VPWR U$$4231/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater548 U$$2542/A2 VGND VGND VPWR VPWR U$$2524/A2 sky130_fd_sc_hd__buf_6
Xrepeater559 U$$2196/X VGND VGND VPWR VPWR U$$2308/A2 sky130_fd_sc_hd__buf_4
XFILLER_65_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4241 U$$4241/A U$$4247/A VGND VGND VPWR VPWR U$$4241/X sky130_fd_sc_hd__xor2_1
XU$$4252 U$$4250/B input58/X input59/X U$$4247/Y VGND VGND VPWR VPWR U$$4252/X sky130_fd_sc_hd__a22o_4
XU$$4263 U$$4400/A1 U$$4381/A2 U$$4402/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4264/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_47_2 dadda_fa_2_47_2/A dadda_fa_2_47_2/B dadda_fa_2_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/A dadda_fa_3_47_3/A sky130_fd_sc_hd__fa_1
XU$$4274 U$$4274/A U$$4294/B VGND VGND VPWR VPWR U$$4274/X sky130_fd_sc_hd__xor2_1
XU$$3540 U$$3540/A U$$3550/B VGND VGND VPWR VPWR U$$3540/X sky130_fd_sc_hd__xor2_1
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4285 input71/X U$$4369/A2 input72/X U$$4369/B2 VGND VGND VPWR VPWR U$$4286/A sky130_fd_sc_hd__a22o_1
XU$$3551 U$$3551/A1 U$$3559/A2 input121/X U$$3559/B2 VGND VGND VPWR VPWR U$$3552/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_24_1 dadda_fa_5_24_1/A dadda_fa_5_24_1/B dadda_fa_5_24_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_25_0/B dadda_fa_7_24_0/A sky130_fd_sc_hd__fa_2
XU$$4296 U$$4296/A U$$4310/B VGND VGND VPWR VPWR U$$4296/X sky130_fd_sc_hd__xor2_1
XFILLER_129_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3562 input47/X VGND VGND VPWR VPWR U$$3562/Y sky130_fd_sc_hd__inv_1
XU$$3573 U$$3573/A U$$3665/B VGND VGND VPWR VPWR U$$3573/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_17_0 dadda_fa_5_17_0/A dadda_fa_5_17_0/B dadda_fa_5_17_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_18_0/A dadda_fa_6_17_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_20_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3584 U$$4269/A1 U$$3612/A2 U$$3584/B1 U$$3612/B2 VGND VGND VPWR VPWR U$$3585/A
+ sky130_fd_sc_hd__a22o_1
XU$$2850 U$$4494/A1 U$$2874/A2 U$$4496/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2851/A
+ sky130_fd_sc_hd__a22o_1
XU$$3595 U$$3595/A U$$3613/B VGND VGND VPWR VPWR U$$3595/X sky130_fd_sc_hd__xor2_1
XFILLER_209_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2861 U$$2861/A U$$2869/B VGND VGND VPWR VPWR U$$2861/X sky130_fd_sc_hd__xor2_1
XFILLER_80_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2872 U$$3555/B1 U$$2874/A2 U$$3557/B1 U$$2874/B2 VGND VGND VPWR VPWR U$$2873/A
+ sky130_fd_sc_hd__a22o_1
XU$$2883 U$$2883/A1 U$$2921/A2 U$$3159/A1 U$$2921/B2 VGND VGND VPWR VPWR U$$2884/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2894 U$$2894/A U$$2922/B VGND VGND VPWR VPWR U$$2894/X sky130_fd_sc_hd__xor2_1
XFILLER_205_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1076 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$801 final_adder.U$$800/B final_adder.U$$721/X final_adder.U$$689/X
+ VGND VGND VPWR VPWR final_adder.U$$801/X sky130_fd_sc_hd__a21o_1
XTAP_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$823 final_adder.U$$790/A final_adder.U$$623/X final_adder.U$$711/X
+ VGND VGND VPWR VPWR final_adder.U$$823/X sky130_fd_sc_hd__a21o_1
XTAP_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$845 final_adder.U$$748/X final_adder.U$$813/X final_adder.U$$749/X
+ VGND VGND VPWR VPWR final_adder.U$$845/X sky130_fd_sc_hd__a21o_2
XFILLER_21_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$867 final_adder.U$$770/X final_adder.U$$723/X final_adder.U$$771/X
+ VGND VGND VPWR VPWR final_adder.U$$867/X sky130_fd_sc_hd__a21o_1
XU$$706 U$$706/A U$$712/B VGND VGND VPWR VPWR U$$706/X sky130_fd_sc_hd__xor2_1
XFILLER_29_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$717 U$$717/A1 U$$739/A2 U$$854/B1 U$$739/B2 VGND VGND VPWR VPWR U$$718/A sky130_fd_sc_hd__a22o_1
XFILLER_205_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$889 final_adder.U$$792/X final_adder.U$$625/X final_adder.U$$793/X
+ VGND VGND VPWR VPWR final_adder.U$$889/X sky130_fd_sc_hd__a21o_1
XU$$728 U$$728/A U$$750/B VGND VGND VPWR VPWR U$$728/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_42_1 U$$490/X U$$623/X U$$756/X VGND VGND VPWR VPWR dadda_fa_2_43_3/B
+ dadda_fa_2_42_5/A sky130_fd_sc_hd__fa_1
XFILLER_72_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$739 U$$52/B1 U$$739/A2 U$$56/A1 U$$739/B2 VGND VGND VPWR VPWR U$$740/A sky130_fd_sc_hd__a22o_1
XFILLER_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1606 U$$2165/A1 VGND VGND VPWR VPWR U$$2711/B1 sky130_fd_sc_hd__buf_4
XFILLER_125_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1617 U$$3944/A1 VGND VGND VPWR VPWR U$$4492/A1 sky130_fd_sc_hd__buf_6
XFILLER_192_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1628 U$$2206/B1 VGND VGND VPWR VPWR U$$1932/B1 sky130_fd_sc_hd__buf_4
Xrepeater1639 U$$517/A1 VGND VGND VPWR VPWR U$$928/A1 sky130_fd_sc_hd__buf_6
XFILLER_193_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_71_3 dadda_fa_3_71_3/A dadda_fa_3_71_3/B dadda_fa_3_71_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_72_1/B dadda_fa_4_71_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_156_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_64_2 dadda_fa_3_64_2/A dadda_fa_3_64_2/B dadda_fa_3_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_1/A dadda_fa_4_64_2/B sky130_fd_sc_hd__fa_1
XFILLER_0_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_57_1 dadda_fa_3_57_1/A dadda_fa_3_57_1/B dadda_fa_3_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_0/CIN dadda_fa_4_57_2/A sky130_fd_sc_hd__fa_1
XFILLER_48_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_34_0 dadda_fa_6_34_0/A dadda_fa_6_34_0/B dadda_fa_6_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_35_0/B dadda_fa_7_34_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2102 U$$2102/A U$$2114/B VGND VGND VPWR VPWR U$$2102/X sky130_fd_sc_hd__xor2_1
XU$$2113 U$$3618/B1 U$$2113/A2 U$$2113/B1 U$$2113/B2 VGND VGND VPWR VPWR U$$2114/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2124 U$$2124/A U$$2150/B VGND VGND VPWR VPWR U$$2124/X sky130_fd_sc_hd__xor2_1
XFILLER_74_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2135 U$$3366/B1 U$$2177/A2 U$$2409/B1 U$$2177/B2 VGND VGND VPWR VPWR U$$2136/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1401 U$$1401/A U$$1405/B VGND VGND VPWR VPWR U$$1401/X sky130_fd_sc_hd__xor2_1
XU$$2146 U$$2146/A U$$2184/B VGND VGND VPWR VPWR U$$2146/X sky130_fd_sc_hd__xor2_1
XU$$1412 U$$864/A1 U$$1434/A2 U$$864/B1 U$$1434/B2 VGND VGND VPWR VPWR U$$1413/A sky130_fd_sc_hd__a22o_1
XFILLER_62_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2157 U$$2292/B1 U$$2189/A2 U$$789/A1 U$$2189/B2 VGND VGND VPWR VPWR U$$2158/A
+ sky130_fd_sc_hd__a22o_1
XU$$1423 U$$1423/A U$$1423/B VGND VGND VPWR VPWR U$$1423/X sky130_fd_sc_hd__xor2_1
XFILLER_50_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2168 U$$2168/A input25/X VGND VGND VPWR VPWR U$$2168/X sky130_fd_sc_hd__xor2_1
XU$$2179 U$$4508/A1 U$$2059/X U$$4510/A1 U$$2060/X VGND VGND VPWR VPWR U$$2180/A sky130_fd_sc_hd__a22o_1
XU$$1434 U$$610/B1 U$$1434/A2 U$$477/A1 U$$1434/B2 VGND VGND VPWR VPWR U$$1435/A sky130_fd_sc_hd__a22o_1
XU$$1445 U$$1445/A U$$1449/B VGND VGND VPWR VPWR U$$1445/X sky130_fd_sc_hd__xor2_1
XU$$1456 U$$2415/A1 U$$1462/A2 U$$2415/B1 U$$1462/B2 VGND VGND VPWR VPWR U$$1457/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3294_1747 VGND VGND VPWR VPWR U$$3294_1747/HI U$$3294/A1 sky130_fd_sc_hd__conb_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1467 U$$1467/A U$$1506/A VGND VGND VPWR VPWR U$$1467/X sky130_fd_sc_hd__xor2_1
XU$$1478 U$$2026/A1 U$$1504/A2 U$$932/A1 U$$1504/B2 VGND VGND VPWR VPWR U$$1479/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1489 U$$1489/A U$$1499/B VGND VGND VPWR VPWR U$$1489/X sky130_fd_sc_hd__xor2_1
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_332 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_754 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_107_0 dadda_fa_7_107_0/A dadda_fa_7_107_0/B dadda_fa_7_107_0/CIN VGND
+ VGND VPWR VPWR _404_/D _275_/D sky130_fd_sc_hd__fa_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$108 _404_/Q _276_/Q VGND VGND VPWR VPWR final_adder.U$$917/B1 final_adder.U$$146/A
+ sky130_fd_sc_hd__ha_1
XFILLER_170_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$119 _415_/Q _287_/Q VGND VGND VPWR VPWR final_adder.U$$137/B1 final_adder.U$$136/B
+ sky130_fd_sc_hd__ha_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_52_0 dadda_fa_2_52_0/A dadda_fa_2_52_0/B dadda_fa_2_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_0/B dadda_fa_3_52_2/B sky130_fd_sc_hd__fa_1
XFILLER_38_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4060 U$$4060/A U$$4078/B VGND VGND VPWR VPWR U$$4060/X sky130_fd_sc_hd__xor2_1
XFILLER_54_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater389 U$$1057/A2 VGND VGND VPWR VPWR U$$965/A2 sky130_fd_sc_hd__buf_6
XU$$4071 input104/X U$$4101/A2 input105/X U$$4101/B2 VGND VGND VPWR VPWR U$$4072/A
+ sky130_fd_sc_hd__a22o_1
XU$$4082 U$$4082/A U$$4100/B VGND VGND VPWR VPWR U$$4082/X sky130_fd_sc_hd__xor2_1
XU$$4093 U$$4365/B1 U$$4103/A2 U$$4095/A1 U$$4103/B2 VGND VGND VPWR VPWR U$$4094/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3370 U$$3644/A1 U$$3374/A2 U$$3644/B1 U$$3374/B2 VGND VGND VPWR VPWR U$$3371/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3381 U$$3381/A U$$3389/B VGND VGND VPWR VPWR U$$3381/X sky130_fd_sc_hd__xor2_1
XU$$3392 U$$3801/B1 U$$3394/A2 U$$4077/B1 U$$3394/B2 VGND VGND VPWR VPWR U$$3393/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_6_0 U$$19/X U$$152/X U$$285/X VGND VGND VPWR VPWR dadda_fa_6_7_0/A dadda_fa_6_6_0/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2680 U$$2680/A U$$2680/B VGND VGND VPWR VPWR U$$2680/X sky130_fd_sc_hd__xor2_1
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2691 U$$2691/A1 U$$2691/A2 U$$4335/B1 U$$2691/B2 VGND VGND VPWR VPWR U$$2692/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1990 U$$2810/B1 U$$1990/A2 U$$483/B1 U$$1990/B2 VGND VGND VPWR VPWR U$$1991/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_81_2 dadda_fa_4_81_2/A dadda_fa_4_81_2/B dadda_fa_4_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_82_0/CIN dadda_fa_5_81_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_74_1 dadda_fa_4_74_1/A dadda_fa_4_74_1/B dadda_fa_4_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/B dadda_fa_5_74_1/B sky130_fd_sc_hd__fa_1
XFILLER_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_51_0 dadda_fa_7_51_0/A dadda_fa_7_51_0/B dadda_fa_7_51_0/CIN VGND VGND
+ VPWR VPWR _348_/D _219_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_67_0 dadda_fa_4_67_0/A dadda_fa_4_67_0/B dadda_fa_4_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/A dadda_fa_5_67_1/A sky130_fd_sc_hd__fa_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput104 b[45] VGND VGND VPWR VPWR input104/X sky130_fd_sc_hd__buf_6
XFILLER_153_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput115 b[55] VGND VGND VPWR VPWR input115/X sky130_fd_sc_hd__buf_6
XFILLER_163_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput126 b[7] VGND VGND VPWR VPWR input126/X sky130_fd_sc_hd__buf_8
XTAP_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput137 c[107] VGND VGND VPWR VPWR input137/X sky130_fd_sc_hd__buf_4
XFILLER_114_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput148 c[117] VGND VGND VPWR VPWR input148/X sky130_fd_sc_hd__clkbuf_4
XTAP_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput159 c[127] VGND VGND VPWR VPWR input159/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$631 final_adder.U$$630/B final_adder.U$$527/X final_adder.U$$511/X
+ VGND VGND VPWR VPWR final_adder.U$$631/X sky130_fd_sc_hd__a21o_1
XTAP_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$642 final_adder.U$$658/B final_adder.U$$642/B VGND VGND VPWR VPWR
+ final_adder.U$$754/B sky130_fd_sc_hd__and2_1
XTAP_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$653 final_adder.U$$652/B final_adder.U$$549/X final_adder.U$$533/X
+ VGND VGND VPWR VPWR final_adder.U$$653/X sky130_fd_sc_hd__a21o_1
XTAP_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$664 final_adder.U$$680/B final_adder.U$$664/B VGND VGND VPWR VPWR
+ final_adder.U$$776/B sky130_fd_sc_hd__and2_1
XTAP_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$503 U$$640/A1 U$$527/A2 U$$916/A1 U$$527/B2 VGND VGND VPWR VPWR U$$504/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$675 final_adder.U$$674/B final_adder.U$$571/X final_adder.U$$555/X
+ VGND VGND VPWR VPWR final_adder.U$$675/X sky130_fd_sc_hd__a21o_1
XU$$514 U$$514/A U$$516/B VGND VGND VPWR VPWR U$$514/X sky130_fd_sc_hd__xor2_1
XTAP_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$686 final_adder.U$$702/B final_adder.U$$686/B VGND VGND VPWR VPWR
+ final_adder.U$$798/B sky130_fd_sc_hd__and2_1
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$525 U$$660/B1 U$$527/A2 U$$527/A1 U$$527/B2 VGND VGND VPWR VPWR U$$526/A sky130_fd_sc_hd__a22o_1
XFILLER_72_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater890 U$$80/B2 VGND VGND VPWR VPWR U$$50/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$697 final_adder.U$$696/B final_adder.U$$593/X final_adder.U$$577/X
+ VGND VGND VPWR VPWR final_adder.U$$697/X sky130_fd_sc_hd__a21o_1
XTAP_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$536 U$$536/A U$$536/B VGND VGND VPWR VPWR U$$536/X sky130_fd_sc_hd__xor2_1
XTAP_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$547 U$$548/A VGND VGND VPWR VPWR U$$547/Y sky130_fd_sc_hd__inv_1
XU$$558 U$$969/A1 U$$578/A2 U$$969/B1 U$$578/B2 VGND VGND VPWR VPWR U$$559/A sky130_fd_sc_hd__a22o_1
XFILLER_147_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$569 U$$569/A U$$579/B VGND VGND VPWR VPWR U$$569/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk _239_/CLK VGND VGND VPWR VPWR _370_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_398 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1403 input25/X VGND VGND VPWR VPWR U$$2184/B sky130_fd_sc_hd__buf_6
XFILLER_197_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1414 U$$2017/B VGND VGND VPWR VPWR U$$1991/B sky130_fd_sc_hd__buf_12
XFILLER_181_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1425 U$$1914/B VGND VGND VPWR VPWR U$$1878/B sky130_fd_sc_hd__buf_12
XFILLER_197_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1436 U$$1780/A VGND VGND VPWR VPWR U$$1765/B sky130_fd_sc_hd__buf_12
XFILLER_158_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1447 U$$1423/B VGND VGND VPWR VPWR U$$1399/B sky130_fd_sc_hd__buf_6
XFILLER_181_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1458 U$$2901/B1 VGND VGND VPWR VPWR U$$2492/A1 sky130_fd_sc_hd__clkbuf_4
Xrepeater1469 input127/X VGND VGND VPWR VPWR U$$24/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_730 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_774 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4387_1768 VGND VGND VPWR VPWR U$$4387_1768/HI U$$4387/A sky130_fd_sc_hd__conb_1
XFILLER_36_947 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1220 U$$944/B1 U$$1222/A2 U$$811/A1 U$$1222/B2 VGND VGND VPWR VPWR U$$1221/A sky130_fd_sc_hd__a22o_1
XU$$1231 U$$1231/A U$$1232/A VGND VGND VPWR VPWR U$$1231/X sky130_fd_sc_hd__xor2_1
XU$$1242 U$$1242/A U$$1272/B VGND VGND VPWR VPWR U$$1242/X sky130_fd_sc_hd__xor2_1
XFILLER_206_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1253 U$$1799/B1 U$$1271/A2 U$$1666/A1 U$$1281/B2 VGND VGND VPWR VPWR U$$1254/A
+ sky130_fd_sc_hd__a22o_1
XU$$1264 U$$1264/A U$$1270/B VGND VGND VPWR VPWR U$$1264/X sky130_fd_sc_hd__xor2_1
XU$$1275 U$$864/A1 U$$1323/A2 U$$864/B1 U$$1307/B2 VGND VGND VPWR VPWR U$$1276/A sky130_fd_sc_hd__a22o_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_42_clk _385_/CLK VGND VGND VPWR VPWR _422_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_188_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1286 U$$1286/A U$$1286/B VGND VGND VPWR VPWR U$$1286/X sky130_fd_sc_hd__xor2_1
XFILLER_149_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1297 U$$3213/B1 U$$1323/A2 U$$477/A1 U$$1349/B2 VGND VGND VPWR VPWR U$$1298/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_91_1 dadda_fa_5_91_1/A dadda_fa_5_91_1/B dadda_fa_5_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_92_0/B dadda_fa_7_91_0/A sky130_fd_sc_hd__fa_1
XFILLER_163_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_84_0 dadda_fa_5_84_0/A dadda_fa_5_84_0/B dadda_fa_5_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_85_0/A dadda_fa_6_84_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_1166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1080 final_adder.U$$198/A final_adder.U$$811/X VGND VGND VPWR VPWR
+ output336/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1091 final_adder.U$$188/B final_adder.U$$959/X VGND VGND VPWR VPWR
+ output348/A sky130_fd_sc_hd__xor2_1
XFILLER_172_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_76_7 U$$4282/X U$$4415/X input230/X VGND VGND VPWR VPWR dadda_fa_2_77_2/CIN
+ dadda_fa_2_76_5/CIN sky130_fd_sc_hd__fa_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_6 dadda_fa_1_69_6/A dadda_fa_1_69_6/B dadda_fa_1_69_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_2/B dadda_fa_2_69_5/B sky130_fd_sc_hd__fa_1
XFILLER_133_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _200_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_33_clk _255_/CLK VGND VGND VPWR VPWR _419_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_99_0 dadda_fa_7_99_0/A dadda_fa_7_99_0/B dadda_fa_7_99_0/CIN VGND VGND
+ VPWR VPWR _396_/D _267_/D sky130_fd_sc_hd__fa_1
XFILLER_33_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4453_1803 VGND VGND VPWR VPWR U$$4453_1803/HI U$$4453/B sky130_fd_sc_hd__conb_1
Xdadda_fa_3_100_2 dadda_fa_3_100_2/A dadda_fa_3_100_2/B dadda_fa_3_100_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_1/A dadda_fa_4_100_2/B sky130_fd_sc_hd__fa_1
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_64_5 U$$2130/X U$$2263/X U$$2396/X VGND VGND VPWR VPWR dadda_fa_1_65_7/A
+ dadda_fa_2_64_0/A sky130_fd_sc_hd__fa_1
XTAP_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_114_0 dadda_fa_6_114_0/A dadda_fa_6_114_0/B dadda_fa_6_114_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_115_0/B dadda_fa_7_114_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$450 final_adder.U$$454/B final_adder.U$$450/B VGND VGND VPWR VPWR
+ final_adder.U$$574/B sky130_fd_sc_hd__and2_1
XTAP_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$300 U$$26/A1 U$$302/A2 U$$28/A1 U$$302/B2 VGND VGND VPWR VPWR U$$301/A sky130_fd_sc_hd__a22o_1
XFILLER_18_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$461 final_adder.U$$460/B final_adder.U$$339/X final_adder.U$$335/X
+ VGND VGND VPWR VPWR final_adder.U$$461/X sky130_fd_sc_hd__a21o_1
XTAP_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$472 final_adder.U$$476/B final_adder.U$$472/B VGND VGND VPWR VPWR
+ final_adder.U$$596/B sky130_fd_sc_hd__and2_1
XTAP_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$311 U$$311/A U$$343/B VGND VGND VPWR VPWR U$$311/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$483 final_adder.U$$482/B final_adder.U$$361/X final_adder.U$$357/X
+ VGND VGND VPWR VPWR final_adder.U$$483/X sky130_fd_sc_hd__a21o_1
XTAP_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$322 U$$733/A1 U$$350/A2 U$$48/B1 U$$350/B2 VGND VGND VPWR VPWR U$$323/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_34_3 dadda_fa_3_34_3/A dadda_fa_3_34_3/B dadda_fa_3_34_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_35_1/B dadda_fa_4_34_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$494 final_adder.U$$498/B final_adder.U$$494/B VGND VGND VPWR VPWR
+ final_adder.U$$610/A sky130_fd_sc_hd__and2_1
XTAP_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$333 U$$333/A U$$351/B VGND VGND VPWR VPWR U$$333/X sky130_fd_sc_hd__xor2_1
XTAP_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$344 U$$70/A1 U$$366/A2 U$$72/A1 U$$366/B2 VGND VGND VPWR VPWR U$$345/A sky130_fd_sc_hd__a22o_1
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_27_2 input176/X dadda_fa_3_27_2/B dadda_fa_3_27_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_28_1/A dadda_fa_4_27_2/B sky130_fd_sc_hd__fa_1
XU$$355 U$$355/A U$$397/B VGND VGND VPWR VPWR U$$355/X sky130_fd_sc_hd__xor2_1
XTAP_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$366 U$$366/A1 U$$366/A2 U$$916/A1 U$$366/B2 VGND VGND VPWR VPWR U$$367/A sky130_fd_sc_hd__a22o_1
XU$$377 U$$377/A U$$377/B VGND VGND VPWR VPWR U$$377/X sky130_fd_sc_hd__xor2_1
XFILLER_72_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$388 U$$660/B1 U$$394/A2 U$$388/B1 U$$394/B2 VGND VGND VPWR VPWR U$$389/A sky130_fd_sc_hd__a22o_1
XFILLER_199_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$399 U$$399/A U$$411/A VGND VGND VPWR VPWR U$$399/X sky130_fd_sc_hd__xor2_1
XFILLER_199_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_24_clk _380_/CLK VGND VGND VPWR VPWR _390_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1200 U$$2609/B1 VGND VGND VPWR VPWR U$$1515/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_148_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1211 U$$673/B VGND VGND VPWR VPWR U$$625/B sky130_fd_sc_hd__buf_6
Xrepeater1222 U$$548/A VGND VGND VPWR VPWR U$$546/B sky130_fd_sc_hd__buf_6
Xrepeater1233 U$$4243/B VGND VGND VPWR VPWR U$$4165/B sky130_fd_sc_hd__buf_6
XFILLER_5_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1244 U$$367/B VGND VGND VPWR VPWR U$$343/B sky130_fd_sc_hd__buf_6
XFILLER_99_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1255 U$$4109/A VGND VGND VPWR VPWR U$$4044/B sky130_fd_sc_hd__buf_8
XFILLER_154_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1266 input53/X VGND VGND VPWR VPWR U$$3971/B sky130_fd_sc_hd__buf_6
Xrepeater1277 U$$958/A VGND VGND VPWR VPWR U$$919/B sky130_fd_sc_hd__buf_6
XFILLER_99_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1288 U$$3697/B VGND VGND VPWR VPWR U$$3683/B sky130_fd_sc_hd__buf_6
XFILLER_10_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1299 U$$3518/B VGND VGND VPWR VPWR U$$3480/B sky130_fd_sc_hd__buf_12
XFILLER_45_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_79_5 dadda_fa_2_79_5/A dadda_fa_2_79_5/B dadda_fa_2_79_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_80_2/A dadda_fa_4_79_0/A sky130_fd_sc_hd__fa_2
XU$$1924_1725 VGND VGND VPWR VPWR U$$1924_1725/HI U$$1924/A1 sky130_fd_sc_hd__conb_1
XFILLER_68_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_30_4 U$$1663/X U$$1796/X VGND VGND VPWR VPWR dadda_fa_3_31_2/B dadda_fa_4_30_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_122_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_7_0_0 U$$7/X U$$9/B VGND VGND VPWR VPWR _297_/D _168_/D sky130_fd_sc_hd__ha_1
XFILLER_36_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_clk _219_/CLK VGND VGND VPWR VPWR _218_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1050 U$$1050/A U$$968/B VGND VGND VPWR VPWR U$$1050/X sky130_fd_sc_hd__xor2_1
XFILLER_211_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1061 U$$924/A1 U$$993/A2 U$$926/A1 U$$993/B2 VGND VGND VPWR VPWR U$$1062/A sky130_fd_sc_hd__a22o_1
XFILLER_204_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1072 U$$1072/A U$$962/A VGND VGND VPWR VPWR U$$1072/X sky130_fd_sc_hd__xor2_1
XFILLER_52_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1083 U$$944/B1 U$$1083/A2 U$$811/A1 U$$1083/B2 VGND VGND VPWR VPWR U$$1084/A sky130_fd_sc_hd__a22o_1
XFILLER_143_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1094 U$$1094/A U$$1095/A VGND VGND VPWR VPWR U$$1094/X sky130_fd_sc_hd__xor2_1
XFILLER_192_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_82_7 U$$4028/X U$$4161/X VGND VGND VPWR VPWR dadda_fa_2_83_3/CIN dadda_fa_3_82_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_192_947 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_109_1 dadda_fa_5_109_1/A dadda_fa_5_109_1/B dadda_fa_5_109_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_110_0/B dadda_fa_7_109_0/A sky130_fd_sc_hd__fa_2
XFILLER_160_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_81_5 U$$3228/X U$$3361/X U$$3494/X VGND VGND VPWR VPWR dadda_fa_2_82_2/CIN
+ dadda_fa_2_81_5/B sky130_fd_sc_hd__fa_1
XFILLER_104_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_74_4 U$$3347/X U$$3480/X U$$3613/X VGND VGND VPWR VPWR dadda_fa_2_75_1/CIN
+ dadda_fa_2_74_4/CIN sky130_fd_sc_hd__fa_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_3 U$$3732/X U$$3865/X U$$3998/X VGND VGND VPWR VPWR dadda_fa_2_68_1/B
+ dadda_fa_2_67_4/B sky130_fd_sc_hd__fa_1
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_44_2 dadda_fa_4_44_2/A dadda_fa_4_44_2/B dadda_fa_4_44_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_45_0/CIN dadda_fa_5_44_1/CIN sky130_fd_sc_hd__fa_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4116_1761 VGND VGND VPWR VPWR U$$4116_1761/HI U$$4116/A1 sky130_fd_sc_hd__conb_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4483_1818 VGND VGND VPWR VPWR U$$4483_1818/HI U$$4483/B sky130_fd_sc_hd__conb_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_37_1 dadda_fa_4_37_1/A dadda_fa_4_37_1/B dadda_fa_4_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/B dadda_fa_5_37_1/B sky130_fd_sc_hd__fa_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_14_0 dadda_fa_7_14_0/A dadda_fa_7_14_0/B dadda_fa_7_14_0/CIN VGND VGND
+ VPWR VPWR _311_/D _182_/D sky130_fd_sc_hd__fa_1
XFILLER_26_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_270_ _399_/CLK _270_/D VGND VGND VPWR VPWR _270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_782 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_62_2 U$$929/X U$$1062/X U$$1195/X VGND VGND VPWR VPWR dadda_fa_1_63_6/A
+ dadda_fa_1_62_8/A sky130_fd_sc_hd__fa_1
XTAP_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3903 U$$3903/A U$$3903/B VGND VGND VPWR VPWR U$$3903/X sky130_fd_sc_hd__xor2_1
XFILLER_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3914 U$$4049/B1 U$$3966/A2 input94/X U$$3966/B2 VGND VGND VPWR VPWR U$$3915/A
+ sky130_fd_sc_hd__a22o_1
XU$$3925 U$$3925/A U$$3927/B VGND VGND VPWR VPWR U$$3925/X sky130_fd_sc_hd__xor2_1
XTAP_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3936 U$$4484/A1 U$$3966/A2 U$$4484/B1 U$$3966/B2 VGND VGND VPWR VPWR U$$3937/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3947 U$$3947/A U$$3947/B VGND VGND VPWR VPWR U$$3947/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_32_0 U$$2227/B input182/X dadda_fa_3_32_0/CIN VGND VGND VPWR VPWR dadda_fa_4_33_0/B
+ dadda_fa_4_32_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$280 final_adder.U$$282/B final_adder.U$$280/B VGND VGND VPWR VPWR
+ final_adder.U$$406/B sky130_fd_sc_hd__and2_1
XTAP_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3958 U$$4095/A1 U$$3968/A2 U$$3960/A1 U$$3968/B2 VGND VGND VPWR VPWR U$$3959/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$291 final_adder.U$$290/B final_adder.U$$165/X final_adder.U$$163/X
+ VGND VGND VPWR VPWR final_adder.U$$291/X sky130_fd_sc_hd__a21o_1
XTAP_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3969 U$$3969/A U$$3972/A VGND VGND VPWR VPWR U$$3969/X sky130_fd_sc_hd__xor2_1
XU$$130 U$$676/B1 U$$4/X U$$678/B1 U$$5/X VGND VGND VPWR VPWR U$$131/A sky130_fd_sc_hd__a22o_1
XTAP_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$141 U$$139/Y U$$138/A U$$3/A U$$140/X U$$137/Y VGND VGND VPWR VPWR U$$141/X sky130_fd_sc_hd__a32o_4
XFILLER_40_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$152 U$$152/A U$$176/B VGND VGND VPWR VPWR U$$152/X sky130_fd_sc_hd__xor2_1
XTAP_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$163 U$$26/A1 U$$165/A2 U$$28/A1 U$$165/B2 VGND VGND VPWR VPWR U$$164/A sky130_fd_sc_hd__a22o_1
XTAP_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$174 U$$174/A U$$176/B VGND VGND VPWR VPWR U$$174/X sky130_fd_sc_hd__xor2_1
XFILLER_33_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$185 U$$48/A1 U$$209/A2 U$$48/B1 U$$209/B2 VGND VGND VPWR VPWR U$$186/A sky130_fd_sc_hd__a22o_1
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$196 U$$196/A U$$218/B VGND VGND VPWR VPWR U$$196/X sky130_fd_sc_hd__xor2_1
XFILLER_60_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_399_ _399_/CLK _399_/D VGND VGND VPWR VPWR _399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_91_4 dadda_fa_2_91_4/A dadda_fa_2_91_4/B dadda_fa_2_91_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_92_1/CIN dadda_fa_3_91_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_57_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1030 U$$4311/A1 VGND VGND VPWR VPWR U$$4309/B1 sky130_fd_sc_hd__buf_6
XFILLER_126_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1041 U$$3483/B1 VGND VGND VPWR VPWR U$$2113/B1 sky130_fd_sc_hd__buf_6
Xrepeater1052 U$$56/B1 VGND VGND VPWR VPWR U$$58/A1 sky130_fd_sc_hd__buf_4
XFILLER_142_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_84_3 dadda_fa_2_84_3/A dadda_fa_2_84_3/B dadda_fa_2_84_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/B dadda_fa_3_84_3/B sky130_fd_sc_hd__fa_1
Xrepeater1063 U$$4029/A1 VGND VGND VPWR VPWR U$$4440/A1 sky130_fd_sc_hd__buf_4
XFILLER_5_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1074 U$$52/A1 VGND VGND VPWR VPWR U$$598/B1 sky130_fd_sc_hd__buf_4
Xrepeater1085 U$$2925/B1 VGND VGND VPWR VPWR U$$598/A1 sky130_fd_sc_hd__buf_6
XFILLER_99_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1096 U$$4293/B1 VGND VGND VPWR VPWR U$$3747/A1 sky130_fd_sc_hd__buf_6
XFILLER_173_1259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_77_2 dadda_fa_2_77_2/A dadda_fa_2_77_2/B dadda_fa_2_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/A dadda_fa_3_77_3/A sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_4_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _304_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_54_1 dadda_fa_5_54_1/A dadda_fa_5_54_1/B dadda_fa_5_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_55_0/B dadda_fa_7_54_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_47_0 dadda_fa_5_47_0/A dadda_fa_5_47_0/B dadda_fa_5_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_48_0/A dadda_fa_6_47_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_110_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_100_1 U$$2867/X U$$3000/X U$$3133/X VGND VGND VPWR VPWR dadda_fa_3_101_1/CIN
+ dadda_fa_3_100_3/A sky130_fd_sc_hd__fa_1
XFILLER_169_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3020_1743 VGND VGND VPWR VPWR U$$3020_1743/HI U$$3020/A1 sky130_fd_sc_hd__conb_1
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$280_1739 VGND VGND VPWR VPWR U$$280_1739/HI U$$280/A1 sky130_fd_sc_hd__conb_1
XFILLER_177_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_121_0 U$$4372/X U$$4505/X input153/X VGND VGND VPWR VPWR dadda_fa_6_122_0/A
+ dadda_fa_6_121_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_165_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_110_0_1865 VGND VGND VPWR VPWR dadda_fa_3_110_0/A dadda_fa_3_110_0_1865/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_78_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_72_1 U$$2412/X U$$2545/X U$$2678/X VGND VGND VPWR VPWR dadda_fa_2_73_0/CIN
+ dadda_fa_2_72_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_65_0 U$$2531/X U$$2664/X U$$2797/X VGND VGND VPWR VPWR dadda_fa_2_66_0/B
+ dadda_fa_2_65_3/B sky130_fd_sc_hd__fa_1
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2509 U$$2509/A U$$2597/B VGND VGND VPWR VPWR U$$2509/X sky130_fd_sc_hd__xor2_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1808 U$$1808/A U$$1832/B VGND VGND VPWR VPWR U$$1808/X sky130_fd_sc_hd__xor2_1
XFILLER_27_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1819 U$$860/A1 U$$1819/A2 U$$860/B1 U$$1819/B2 VGND VGND VPWR VPWR U$$1820/A sky130_fd_sc_hd__a22o_1
XFILLER_15_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_322_ _323_/CLK _322_/D VGND VGND VPWR VPWR _322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_253_ _385_/CLK _253_/D VGND VGND VPWR VPWR _253_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_211_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_184_ _337_/CLK _184_/D VGND VGND VPWR VPWR _184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_94_2 dadda_fa_3_94_2/A dadda_fa_3_94_2/B dadda_fa_3_94_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_1/A dadda_fa_4_94_2/B sky130_fd_sc_hd__fa_1
XFILLER_6_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_87_1 dadda_fa_3_87_1/A dadda_fa_3_87_1/B dadda_fa_3_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_0/CIN dadda_fa_4_87_2/A sky130_fd_sc_hd__fa_1
XFILLER_163_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_64_0 dadda_fa_6_64_0/A dadda_fa_6_64_0/B dadda_fa_6_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_65_0/B dadda_fa_7_64_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_9_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater708 U$$3968/B2 VGND VGND VPWR VPWR U$$3966/B2 sky130_fd_sc_hd__buf_8
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater719 U$$3644/B2 VGND VGND VPWR VPWR U$$3612/B2 sky130_fd_sc_hd__buf_4
XU$$4401 U$$4401/A U$$4401/B VGND VGND VPWR VPWR U$$4401/X sky130_fd_sc_hd__xor2_1
XFILLER_65_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4412 input66/X U$$4388/X input67/X U$$4426/B2 VGND VGND VPWR VPWR U$$4413/A sky130_fd_sc_hd__a22o_1
XU$$4423 U$$4423/A U$$4423/B VGND VGND VPWR VPWR U$$4423/X sky130_fd_sc_hd__xor2_1
XU$$4434 U$$4434/A1 U$$4388/X U$$4436/A1 U$$4389/X VGND VGND VPWR VPWR U$$4435/A sky130_fd_sc_hd__a22o_1
XFILLER_64_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3700 input50/X VGND VGND VPWR VPWR U$$3702/B sky130_fd_sc_hd__inv_1
XU$$4445 U$$4445/A U$$4445/B VGND VGND VPWR VPWR U$$4445/X sky130_fd_sc_hd__xor2_1
XU$$4456 U$$4456/A1 U$$4388/X U$$4458/A1 U$$4476/B2 VGND VGND VPWR VPWR U$$4457/A
+ sky130_fd_sc_hd__a22o_1
XU$$3711 U$$3846/B1 U$$3753/A2 U$$3713/A1 U$$3753/B2 VGND VGND VPWR VPWR U$$3712/A
+ sky130_fd_sc_hd__a22o_1
XU$$4467 U$$4467/A U$$4467/B VGND VGND VPWR VPWR U$$4467/X sky130_fd_sc_hd__xor2_1
XTAP_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_116_1 U$$4229/X U$$4362/X U$$4495/X VGND VGND VPWR VPWR dadda_fa_5_117_0/B
+ dadda_fa_5_116_1/B sky130_fd_sc_hd__fa_1
XU$$3722 U$$3722/A U$$3740/B VGND VGND VPWR VPWR U$$3722/X sky130_fd_sc_hd__xor2_1
XFILLER_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4478 U$$4478/A1 U$$4388/X U$$4478/B1 U$$4486/B2 VGND VGND VPWR VPWR U$$4479/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3733 U$$4418/A1 U$$3773/A2 U$$4420/A1 U$$3773/B2 VGND VGND VPWR VPWR U$$3734/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3744 U$$3744/A U$$3778/B VGND VGND VPWR VPWR U$$3744/X sky130_fd_sc_hd__xor2_1
XU$$4489 U$$4489/A U$$4489/B VGND VGND VPWR VPWR U$$4489/X sky130_fd_sc_hd__xor2_1
XTAP_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_109_0 dadda_fa_4_109_0/A dadda_fa_4_109_0/B dadda_fa_4_109_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/A dadda_fa_5_109_1/A sky130_fd_sc_hd__fa_1
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3755 U$$4029/A1 U$$3777/A2 input82/X U$$3777/B2 VGND VGND VPWR VPWR U$$3756/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3766 U$$3766/A U$$3774/B VGND VGND VPWR VPWR U$$3766/X sky130_fd_sc_hd__xor2_1
XU$$3777 U$$4049/B1 U$$3777/A2 input94/X U$$3777/B2 VGND VGND VPWR VPWR U$$3778/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3788 U$$3788/A U$$3794/B VGND VGND VPWR VPWR U$$3788/X sky130_fd_sc_hd__xor2_1
XTAP_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3799 U$$4210/A1 U$$3813/A2 U$$4210/B1 U$$3813/B2 VGND VGND VPWR VPWR U$$3800/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_991 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_82_0 U$$4294/X U$$4427/X input237/X VGND VGND VPWR VPWR dadda_fa_3_83_0/B
+ dadda_fa_3_82_2/B sky130_fd_sc_hd__fa_1
XFILLER_114_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_51_6 U$$2503/X U$$2636/X U$$2769/X VGND VGND VPWR VPWR dadda_fa_2_52_2/B
+ dadda_fa_2_51_5/B sky130_fd_sc_hd__fa_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_3_0 input190/X dadda_fa_7_3_0/B dadda_ha_6_3_0/SUM VGND VGND VPWR VPWR
+ _300_/D _171_/D sky130_fd_sc_hd__fa_1
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_81_0 dadda_fa_7_81_0/A dadda_fa_7_81_0/B dadda_fa_7_81_0/CIN VGND VGND
+ VPWR VPWR _378_/D _249_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_97_0 dadda_fa_4_97_0/A dadda_fa_4_97_0/B dadda_fa_4_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/A dadda_fa_5_97_1/A sky130_fd_sc_hd__fa_1
XFILLER_137_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3007 input122/X U$$3011/A2 U$$3555/B1 U$$3011/B2 VGND VGND VPWR VPWR U$$3008/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3018 U$$3016/Y input39/X input38/X U$$3017/X U$$3014/Y VGND VGND VPWR VPWR U$$3018/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3029 U$$3029/A U$$3075/B VGND VGND VPWR VPWR U$$3029/X sky130_fd_sc_hd__xor2_1
XU$$2306 U$$936/A1 U$$2196/X U$$936/B1 U$$2197/X VGND VGND VPWR VPWR U$$2307/A sky130_fd_sc_hd__a22o_1
XFILLER_74_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2317 U$$2317/A U$$2317/B VGND VGND VPWR VPWR U$$2317/X sky130_fd_sc_hd__xor2_1
XU$$2328 U$$2328/A VGND VGND VPWR VPWR U$$2328/Y sky130_fd_sc_hd__inv_1
XFILLER_76_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2339 U$$3296/B1 U$$2417/A2 U$$3300/A1 U$$2417/B2 VGND VGND VPWR VPWR U$$2340/A
+ sky130_fd_sc_hd__a22o_1
XU$$1605 U$$2016/A1 U$$1607/A2 U$$2975/B1 U$$1607/B2 VGND VGND VPWR VPWR U$$1606/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1616 U$$1616/A U$$1628/B VGND VGND VPWR VPWR U$$1616/X sky130_fd_sc_hd__xor2_1
XFILLER_15_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1627 U$$2449/A1 U$$1635/A2 U$$1764/B1 U$$1635/B2 VGND VGND VPWR VPWR U$$1628/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1638 U$$1638/A U$$1638/B VGND VGND VPWR VPWR U$$1638/X sky130_fd_sc_hd__xor2_1
XU$$1649 U$$1647/B input16/X input17/X U$$1644/Y VGND VGND VPWR VPWR U$$1649/X sky130_fd_sc_hd__a22o_2
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_76 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_305_ _326_/CLK _305_/D VGND VGND VPWR VPWR _305_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_236_ _367_/CLK _236_/D VGND VGND VPWR VPWR _236_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_155_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_61_5 dadda_fa_2_61_5/A dadda_fa_2_61_5/B dadda_fa_2_61_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_62_2/A dadda_fa_4_61_0/A sky130_fd_sc_hd__fa_2
Xrepeater505 U$$3018/X VGND VGND VPWR VPWR U$$3098/A2 sky130_fd_sc_hd__buf_6
Xrepeater516 U$$2977/A2 VGND VGND VPWR VPWR U$$2967/A2 sky130_fd_sc_hd__buf_12
XFILLER_111_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater527 U$$2796/A2 VGND VGND VPWR VPWR U$$2790/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_54_4 dadda_fa_2_54_4/A dadda_fa_2_54_4/B dadda_fa_2_54_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_1/CIN dadda_fa_3_54_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater538 U$$2691/A2 VGND VGND VPWR VPWR U$$2683/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4220 U$$4494/A1 U$$4240/A2 input112/X U$$4240/B2 VGND VGND VPWR VPWR U$$4221/A
+ sky130_fd_sc_hd__a22o_1
XU$$4231 U$$4231/A U$$4247/A VGND VGND VPWR VPWR U$$4231/X sky130_fd_sc_hd__xor2_1
XFILLER_1_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater549 U$$2558/A2 VGND VGND VPWR VPWR U$$2542/A2 sky130_fd_sc_hd__buf_8
XFILLER_65_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4242 U$$4379/A1 U$$4114/X U$$4242/B1 U$$4115/X VGND VGND VPWR VPWR U$$4243/A sky130_fd_sc_hd__a22o_1
XU$$4253 U$$4253/A1 U$$4275/A2 U$$4392/A1 U$$4275/B2 VGND VGND VPWR VPWR U$$4254/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_47_3 dadda_fa_2_47_3/A dadda_fa_2_47_3/B dadda_fa_2_47_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/B dadda_fa_3_47_3/B sky130_fd_sc_hd__fa_1
XFILLER_93_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4264 U$$4264/A U$$4384/A VGND VGND VPWR VPWR U$$4264/X sky130_fd_sc_hd__xor2_1
XU$$3530 U$$3530/A U$$3550/B VGND VGND VPWR VPWR U$$3530/X sky130_fd_sc_hd__xor2_1
XFILLER_65_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4275 U$$4275/A1 U$$4275/A2 U$$4275/B1 U$$4275/B2 VGND VGND VPWR VPWR U$$4276/A
+ sky130_fd_sc_hd__a22o_1
XU$$3541 input114/X U$$3559/A2 U$$3817/A1 U$$3559/B2 VGND VGND VPWR VPWR U$$3542/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4286 U$$4286/A U$$4370/B VGND VGND VPWR VPWR U$$4286/X sky130_fd_sc_hd__xor2_1
XU$$3552 U$$3552/A U$$3561/A VGND VGND VPWR VPWR U$$3552/X sky130_fd_sc_hd__xor2_1
XU$$4297 U$$4434/A1 U$$4297/A2 U$$4297/B1 U$$4297/B2 VGND VGND VPWR VPWR U$$4298/A
+ sky130_fd_sc_hd__a22o_1
XU$$3563 input48/X VGND VGND VPWR VPWR U$$3565/B sky130_fd_sc_hd__inv_1
XFILLER_93_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3574 U$$3846/B1 U$$3660/A2 U$$3713/A1 U$$3660/B2 VGND VGND VPWR VPWR U$$3575/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_17_1 dadda_fa_5_17_1/A dadda_fa_5_17_1/B dadda_fa_5_17_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_18_0/B dadda_fa_7_17_0/A sky130_fd_sc_hd__fa_1
XU$$2840 U$$2975/B1 U$$2744/X U$$2842/A1 U$$2745/X VGND VGND VPWR VPWR U$$2841/A sky130_fd_sc_hd__a22o_1
XU$$3585 U$$3585/A U$$3609/B VGND VGND VPWR VPWR U$$3585/X sky130_fd_sc_hd__xor2_1
XU$$2851 U$$2851/A U$$2876/A VGND VGND VPWR VPWR U$$2851/X sky130_fd_sc_hd__xor2_1
XU$$3596 U$$4418/A1 U$$3636/A2 U$$4420/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3597/A
+ sky130_fd_sc_hd__a22o_1
XU$$2862 U$$3684/A1 U$$2868/A2 U$$3547/B1 U$$2868/B2 VGND VGND VPWR VPWR U$$2863/A
+ sky130_fd_sc_hd__a22o_1
XU$$2873 U$$2873/A U$$2876/A VGND VGND VPWR VPWR U$$2873/X sky130_fd_sc_hd__xor2_1
XFILLER_178_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2884 U$$2884/A U$$2922/B VGND VGND VPWR VPWR U$$2884/X sky130_fd_sc_hd__xor2_1
XFILLER_90_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2895 U$$3852/B1 U$$2921/A2 U$$3719/A1 U$$2921/B2 VGND VGND VPWR VPWR U$$2896/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_390 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_755 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_4_120_1 U$$4237/X U$$4370/X VGND VGND VPWR VPWR dadda_fa_5_121_1/B dadda_ha_4_120_1/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_780 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_43_4 U$$1689/X U$$1822/X VGND VGND VPWR VPWR dadda_fa_2_44_4/A dadda_fa_3_43_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$813 final_adder.U$$780/A final_adder.U$$733/X final_adder.U$$701/X
+ VGND VGND VPWR VPWR final_adder.U$$813/X sky130_fd_sc_hd__a21o_1
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_4_13_2 U$$831/X input161/X VGND VGND VPWR VPWR dadda_fa_5_14_0/CIN dadda_ha_4_13_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_60_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$857 final_adder.U$$760/X final_adder.U$$825/X final_adder.U$$761/X
+ VGND VGND VPWR VPWR final_adder.U$$857/X sky130_fd_sc_hd__a21o_2
XFILLER_60_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$707 U$$22/A1 U$$739/A2 U$$983/A1 U$$739/B2 VGND VGND VPWR VPWR U$$708/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$879 final_adder.U$$782/X final_adder.U$$735/X final_adder.U$$783/X
+ VGND VGND VPWR VPWR final_adder.U$$879/X sky130_fd_sc_hd__a21o_2
XU$$718 U$$718/A U$$740/B VGND VGND VPWR VPWR U$$718/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_42_2 U$$889/X U$$1022/X U$$1155/X VGND VGND VPWR VPWR dadda_fa_2_43_3/CIN
+ dadda_fa_2_42_5/B sky130_fd_sc_hd__fa_1
XU$$729 U$$864/B1 U$$749/A2 U$$731/A1 U$$749/B2 VGND VGND VPWR VPWR U$$730/A sky130_fd_sc_hd__a22o_1
XFILLER_186_1236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_12_0 U$$31/X U$$164/X U$$297/X VGND VGND VPWR VPWR dadda_fa_5_13_0/A dadda_fa_5_12_1/A
+ sky130_fd_sc_hd__fa_1
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1607 U$$2165/A1 VGND VGND VPWR VPWR U$$930/B1 sky130_fd_sc_hd__buf_6
Xrepeater1618 input110/X VGND VGND VPWR VPWR U$$3944/A1 sky130_fd_sc_hd__buf_4
Xrepeater1629 U$$975/A1 VGND VGND VPWR VPWR U$$16/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_64_3 dadda_fa_3_64_3/A dadda_fa_3_64_3/B dadda_fa_3_64_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_65_1/B dadda_fa_4_64_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_57_2 dadda_fa_3_57_2/A dadda_fa_3_57_2/B dadda_fa_3_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_1/A dadda_fa_4_57_2/B sky130_fd_sc_hd__fa_1
XFILLER_94_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_891 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_27_0 dadda_fa_6_27_0/A dadda_fa_6_27_0/B dadda_fa_6_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_28_0/B dadda_fa_7_27_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2103 U$$3882/B1 U$$2113/A2 U$$3749/A1 U$$2113/B2 VGND VGND VPWR VPWR U$$2104/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2114 U$$2114/A U$$2114/B VGND VGND VPWR VPWR U$$2114/X sky130_fd_sc_hd__xor2_1
XFILLER_16_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2125 U$$892/A1 U$$2169/A2 U$$894/A1 U$$2169/B2 VGND VGND VPWR VPWR U$$2126/A sky130_fd_sc_hd__a22o_1
XU$$2136 U$$2136/A U$$2178/B VGND VGND VPWR VPWR U$$2136/X sky130_fd_sc_hd__xor2_1
XFILLER_74_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2147 U$$366/A1 U$$2183/A2 U$$2834/A1 U$$2183/B2 VGND VGND VPWR VPWR U$$2148/A
+ sky130_fd_sc_hd__a22o_1
XU$$1402 U$$854/A1 U$$1404/A2 U$$854/B1 U$$1404/B2 VGND VGND VPWR VPWR U$$1403/A sky130_fd_sc_hd__a22o_1
XFILLER_204_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2158 U$$2158/A U$$2191/A VGND VGND VPWR VPWR U$$2158/X sky130_fd_sc_hd__xor2_1
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1413 U$$1413/A U$$1423/B VGND VGND VPWR VPWR U$$1413/X sky130_fd_sc_hd__xor2_1
XFILLER_204_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1424 U$$328/A1 U$$1470/A2 U$$328/B1 U$$1470/B2 VGND VGND VPWR VPWR U$$1425/A sky130_fd_sc_hd__a22o_1
XU$$2169 U$$936/A1 U$$2169/A2 U$$936/B1 U$$2169/B2 VGND VGND VPWR VPWR U$$2170/A sky130_fd_sc_hd__a22o_1
XFILLER_43_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1435 U$$1435/A U$$1459/B VGND VGND VPWR VPWR U$$1435/X sky130_fd_sc_hd__xor2_1
XU$$1446 U$$1446/A1 U$$1448/A2 U$$1448/A1 U$$1448/B2 VGND VGND VPWR VPWR U$$1447/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1457 U$$1457/A U$$1501/B VGND VGND VPWR VPWR U$$1457/X sky130_fd_sc_hd__xor2_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1468 U$$2975/A1 U$$1470/A2 U$$2975/B1 U$$1470/B2 VGND VGND VPWR VPWR U$$1469/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1479 U$$1479/A U$$1501/B VGND VGND VPWR VPWR U$$1479/X sky130_fd_sc_hd__xor2_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_219_ _219_/CLK _219_/D VGND VGND VPWR VPWR _219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$109 _405_/Q _277_/Q VGND VGND VPWR VPWR final_adder.U$$147/B1 final_adder.U$$146/B
+ sky130_fd_sc_hd__ha_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_52_1 dadda_fa_2_52_1/A dadda_fa_2_52_1/B dadda_fa_2_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_0/CIN dadda_fa_3_52_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4050 U$$4050/A U$$4080/B VGND VGND VPWR VPWR U$$4050/X sky130_fd_sc_hd__xor2_1
XU$$4061 U$$4333/B1 U$$4077/A2 U$$912/A1 U$$4077/B2 VGND VGND VPWR VPWR U$$4062/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_45_0 U$$2358/X U$$2491/X U$$2624/X VGND VGND VPWR VPWR dadda_fa_3_46_0/B
+ dadda_fa_3_45_2/B sky130_fd_sc_hd__fa_1
XU$$4072 U$$4072/A U$$4110/A VGND VGND VPWR VPWR U$$4072/X sky130_fd_sc_hd__xor2_1
XFILLER_38_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4083 input111/X U$$4101/A2 input112/X U$$4101/B2 VGND VGND VPWR VPWR U$$4084/A
+ sky130_fd_sc_hd__a22o_1
XU$$4094 U$$4094/A U$$4100/B VGND VGND VPWR VPWR U$$4094/X sky130_fd_sc_hd__xor2_1
XU$$3360 U$$4045/A1 U$$3378/A2 U$$3908/B1 U$$3378/B2 VGND VGND VPWR VPWR U$$3361/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3371 U$$3371/A U$$3375/B VGND VGND VPWR VPWR U$$3371/X sky130_fd_sc_hd__xor2_1
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3382 input102/X U$$3416/A2 input103/X U$$3416/B2 VGND VGND VPWR VPWR U$$3383/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3393 U$$3393/A U$$3395/B VGND VGND VPWR VPWR U$$3393/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2670 U$$2670/A U$$2680/B VGND VGND VPWR VPWR U$$2670/X sky130_fd_sc_hd__xor2_1
XFILLER_62_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2681 U$$4323/B1 U$$2683/A2 U$$4188/B1 U$$2683/B2 VGND VGND VPWR VPWR U$$2682/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2692 U$$2692/A U$$2716/B VGND VGND VPWR VPWR U$$2692/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1980 U$$3348/B1 U$$2016/A2 U$$3215/A1 U$$2016/B2 VGND VGND VPWR VPWR U$$1981/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1991 U$$1991/A U$$1991/B VGND VGND VPWR VPWR U$$1991/X sky130_fd_sc_hd__xor2_1
XFILLER_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_74_2 dadda_fa_4_74_2/A dadda_fa_4_74_2/B dadda_fa_4_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_75_0/CIN dadda_fa_5_74_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_67_1 dadda_fa_4_67_1/A dadda_fa_4_67_1/B dadda_fa_4_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/B dadda_fa_5_67_1/B sky130_fd_sc_hd__fa_1
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput105 b[46] VGND VGND VPWR VPWR input105/X sky130_fd_sc_hd__buf_6
Xinput116 b[56] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__buf_6
XFILLER_130_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_44_0 dadda_fa_7_44_0/A dadda_fa_7_44_0/B dadda_fa_7_44_0/CIN VGND VGND
+ VPWR VPWR _341_/D _212_/D sky130_fd_sc_hd__fa_2
XFILLER_89_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput127 b[8] VGND VGND VPWR VPWR input127/X sky130_fd_sc_hd__buf_12
XTAP_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput138 c[108] VGND VGND VPWR VPWR input138/X sky130_fd_sc_hd__buf_4
XFILLER_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_1_34_0 U$$75/X U$$208/X VGND VGND VPWR VPWR dadda_fa_2_35_5/CIN dadda_fa_3_34_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput149 c[118] VGND VGND VPWR VPWR input149/X sky130_fd_sc_hd__buf_2
XFILLER_57_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$610 final_adder.U$$610/A final_adder.U$$610/B VGND VGND VPWR VPWR
+ final_adder.U$$714/A sky130_fd_sc_hd__and2_1
XTAP_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$621 final_adder.U$$612/A final_adder.U$$505/X final_adder.U$$497/X
+ VGND VGND VPWR VPWR final_adder.U$$621/X sky130_fd_sc_hd__a21o_2
XTAP_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$632 final_adder.U$$648/B final_adder.U$$632/B VGND VGND VPWR VPWR
+ final_adder.U$$744/B sky130_fd_sc_hd__and2_1
XTAP_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$643 final_adder.U$$642/B final_adder.U$$539/X final_adder.U$$523/X
+ VGND VGND VPWR VPWR final_adder.U$$643/X sky130_fd_sc_hd__a21o_1
XTAP_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$654 final_adder.U$$670/B final_adder.U$$654/B VGND VGND VPWR VPWR
+ final_adder.U$$766/B sky130_fd_sc_hd__and2_1
XTAP_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$665 final_adder.U$$664/B final_adder.U$$561/X final_adder.U$$545/X
+ VGND VGND VPWR VPWR final_adder.U$$665/X sky130_fd_sc_hd__a21o_1
XTAP_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$504 U$$504/A U$$504/B VGND VGND VPWR VPWR U$$504/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$676 final_adder.U$$692/B final_adder.U$$676/B VGND VGND VPWR VPWR
+ final_adder.U$$788/B sky130_fd_sc_hd__and2_1
XTAP_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$515 U$$652/A1 U$$515/A2 U$$654/A1 U$$515/B2 VGND VGND VPWR VPWR U$$516/A sky130_fd_sc_hd__a22o_1
Xrepeater880 U$$1174/B2 VGND VGND VPWR VPWR U$$1138/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$687 final_adder.U$$686/B final_adder.U$$583/X final_adder.U$$567/X
+ VGND VGND VPWR VPWR final_adder.U$$687/X sky130_fd_sc_hd__a21o_1
XTAP_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$526 U$$526/A U$$528/B VGND VGND VPWR VPWR U$$526/X sky130_fd_sc_hd__xor2_1
Xrepeater891 U$$134/B2 VGND VGND VPWR VPWR U$$80/B2 sky130_fd_sc_hd__buf_4
XFILLER_99_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$698 final_adder.U$$714/B final_adder.U$$698/B VGND VGND VPWR VPWR
+ final_adder.U$$778/A sky130_fd_sc_hd__and2_1
XTAP_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$537 U$$674/A1 U$$537/A2 U$$676/A1 U$$537/B2 VGND VGND VPWR VPWR U$$538/A sky130_fd_sc_hd__a22o_1
XU$$548 U$$548/A VGND VGND VPWR VPWR U$$548/Y sky130_fd_sc_hd__inv_1
XFILLER_205_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$559 U$$559/A U$$579/B VGND VGND VPWR VPWR U$$559/X sky130_fd_sc_hd__xor2_1
XFILLER_186_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1404 U$$2092/B VGND VGND VPWR VPWR U$$2094/B sky130_fd_sc_hd__buf_6
XFILLER_158_1113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1415 U$$2037/B VGND VGND VPWR VPWR U$$2017/B sky130_fd_sc_hd__buf_8
XFILLER_197_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1426 U$$1914/B VGND VGND VPWR VPWR U$$1917/A sky130_fd_sc_hd__buf_12
Xrepeater1437 input18/X VGND VGND VPWR VPWR U$$1780/A sky130_fd_sc_hd__buf_8
XFILLER_21_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1448 U$$1459/B VGND VGND VPWR VPWR U$$1423/B sky130_fd_sc_hd__buf_6
XFILLER_10_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1459 U$$2901/B1 VGND VGND VPWR VPWR U$$983/B1 sky130_fd_sc_hd__buf_4
XFILLER_180_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_62_0 dadda_fa_3_62_0/A dadda_fa_3_62_0/B dadda_fa_3_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_0/B dadda_fa_4_62_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_786 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_4_9_0 U$$25/X U$$158/X VGND VGND VPWR VPWR dadda_fa_5_10_1/A dadda_ha_4_9_0/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_165_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1210 U$$799/A1 U$$1230/A2 U$$938/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1211/A sky130_fd_sc_hd__a22o_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1221 U$$1221/A U$$1223/B VGND VGND VPWR VPWR U$$1221/X sky130_fd_sc_hd__xor2_1
XFILLER_62_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1232 U$$1232/A VGND VGND VPWR VPWR U$$1232/Y sky130_fd_sc_hd__inv_1
XU$$1243 U$$2202/A1 U$$1311/A2 U$$2202/B1 U$$1271/B2 VGND VGND VPWR VPWR U$$1244/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1254 U$$1254/A U$$1270/B VGND VGND VPWR VPWR U$$1254/X sky130_fd_sc_hd__xor2_1
XFILLER_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1265 U$$854/A1 U$$1271/A2 U$$854/B1 U$$1281/B2 VGND VGND VPWR VPWR U$$1266/A sky130_fd_sc_hd__a22o_1
XFILLER_149_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1276 U$$1276/A U$$1286/B VGND VGND VPWR VPWR U$$1276/X sky130_fd_sc_hd__xor2_1
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1287 U$$328/A1 U$$1337/A2 U$$328/B1 U$$1291/B2 VGND VGND VPWR VPWR U$$1288/A sky130_fd_sc_hd__a22o_1
XU$$1298 U$$1298/A U$$1354/B VGND VGND VPWR VPWR U$$1298/X sky130_fd_sc_hd__xor2_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_84_1 dadda_fa_5_84_1/A dadda_fa_5_84_1/B dadda_fa_5_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_85_0/B dadda_fa_7_84_0/A sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$1070 final_adder.U$$208/A final_adder.U$$821/X VGND VGND VPWR VPWR
+ output325/A sky130_fd_sc_hd__xor2_1
XFILLER_102_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1081 final_adder.U$$198/B final_adder.U$$969/X VGND VGND VPWR VPWR
+ output337/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1092 final_adder.U$$186/A final_adder.U$$895/X VGND VGND VPWR VPWR
+ output349/A sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_77_0 dadda_fa_5_77_0/A dadda_fa_5_77_0/B dadda_fa_5_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_78_0/A dadda_fa_6_77_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_76_8 dadda_fa_1_76_8/A dadda_fa_1_76_8/B dadda_fa_1_76_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_77_3/A dadda_fa_3_76_0/A sky130_fd_sc_hd__fa_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_7 dadda_fa_1_69_7/A dadda_fa_1_69_7/B dadda_fa_1_69_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_2/CIN dadda_fa_2_69_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3190 U$$3190/A U$$3208/B VGND VGND VPWR VPWR U$$3190/X sky130_fd_sc_hd__xor2_1
XFILLER_53_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_100_3 dadda_fa_3_100_3/A dadda_fa_3_100_3/B dadda_fa_3_100_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_101_1/B dadda_fa_4_100_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_95_0 U$$2191/Y U$$2325/X U$$2458/X VGND VGND VPWR VPWR dadda_fa_2_96_5/CIN
+ dadda_fa_3_95_0/A sky130_fd_sc_hd__fa_1
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_474 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_2_108_0 dadda_ha_2_108_0/A U$$3149/X VGND VGND VPWR VPWR dadda_fa_4_109_0/A
+ dadda_fa_4_108_0/A sky130_fd_sc_hd__ha_1
XTAP_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_68_0_1847 VGND VGND VPWR VPWR dadda_fa_0_68_0/A dadda_fa_0_68_0_1847/LO
+ sky130_fd_sc_hd__conb_1
Xfinal_adder.U$$440 final_adder.U$$444/B final_adder.U$$440/B VGND VGND VPWR VPWR
+ final_adder.U$$564/B sky130_fd_sc_hd__and2_1
XTAP_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$451 final_adder.U$$450/B final_adder.U$$329/X final_adder.U$$325/X
+ VGND VGND VPWR VPWR final_adder.U$$451/X sky130_fd_sc_hd__a21o_1
XTAP_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_107_0 dadda_fa_6_107_0/A dadda_fa_6_107_0/B dadda_fa_6_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_108_0/B dadda_fa_7_107_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$462 final_adder.U$$466/B final_adder.U$$462/B VGND VGND VPWR VPWR
+ final_adder.U$$586/B sky130_fd_sc_hd__and2_1
XTAP_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$301 U$$301/A U$$379/B VGND VGND VPWR VPWR U$$301/X sky130_fd_sc_hd__xor2_1
XTAP_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$473 final_adder.U$$472/B final_adder.U$$351/X final_adder.U$$347/X
+ VGND VGND VPWR VPWR final_adder.U$$473/X sky130_fd_sc_hd__a21o_1
XTAP_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$312 U$$312/A1 U$$340/A2 U$$999/A1 U$$340/B2 VGND VGND VPWR VPWR U$$313/A sky130_fd_sc_hd__a22o_1
XTAP_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$484 final_adder.U$$488/B final_adder.U$$484/B VGND VGND VPWR VPWR
+ final_adder.U$$608/B sky130_fd_sc_hd__and2_1
XTAP_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$323 U$$323/A U$$351/B VGND VGND VPWR VPWR U$$323/X sky130_fd_sc_hd__xor2_1
XFILLER_72_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$495 final_adder.U$$494/B final_adder.U$$373/X final_adder.U$$369/X
+ VGND VGND VPWR VPWR final_adder.U$$495/X sky130_fd_sc_hd__a21o_1
XTAP_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$334 U$$745/A1 U$$366/A2 U$$882/B1 U$$366/B2 VGND VGND VPWR VPWR U$$335/A sky130_fd_sc_hd__a22o_1
XTAP_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$345 U$$345/A U$$367/B VGND VGND VPWR VPWR U$$345/X sky130_fd_sc_hd__xor2_1
XFILLER_205_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$356 U$$630/A1 U$$396/A2 U$$630/B1 U$$396/B2 VGND VGND VPWR VPWR U$$357/A sky130_fd_sc_hd__a22o_1
XTAP_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_27_3 dadda_fa_3_27_3/A dadda_fa_3_27_3/B dadda_fa_3_27_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_28_1/B dadda_fa_4_27_2/CIN sky130_fd_sc_hd__fa_1
XU$$367 U$$367/A U$$367/B VGND VGND VPWR VPWR U$$367/X sky130_fd_sc_hd__xor2_1
XFILLER_205_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$378 U$$652/A1 U$$378/A2 U$$654/A1 U$$378/B2 VGND VGND VPWR VPWR U$$379/A sky130_fd_sc_hd__a22o_1
XFILLER_26_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$389 U$$389/A U$$395/B VGND VGND VPWR VPWR U$$389/X sky130_fd_sc_hd__xor2_1
XFILLER_38_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4501_1827 VGND VGND VPWR VPWR U$$4501_1827/HI U$$4501/B sky130_fd_sc_hd__conb_1
XFILLER_199_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_94_0 dadda_fa_6_94_0/A dadda_fa_6_94_0/B dadda_fa_6_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_95_0/B dadda_fa_7_94_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_9_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1201 U$$2609/B1 VGND VGND VPWR VPWR U$$3159/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1212 U$$685/A VGND VGND VPWR VPWR U$$673/B sky130_fd_sc_hd__buf_6
XFILLER_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1223 U$$4294/B VGND VGND VPWR VPWR U$$4278/B sky130_fd_sc_hd__buf_6
XFILLER_181_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1234 U$$4243/B VGND VGND VPWR VPWR U$$4246/A sky130_fd_sc_hd__buf_8
Xrepeater1245 U$$377/B VGND VGND VPWR VPWR U$$379/B sky130_fd_sc_hd__buf_6
XFILLER_99_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1256 input55/X VGND VGND VPWR VPWR U$$4109/A sky130_fd_sc_hd__buf_6
XU$$4393_1773 VGND VGND VPWR VPWR U$$4393_1773/HI U$$4393/B sky130_fd_sc_hd__conb_1
Xrepeater1267 U$$3754/B VGND VGND VPWR VPWR U$$3794/B sky130_fd_sc_hd__buf_6
XFILLER_141_525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1278 U$$945/B VGND VGND VPWR VPWR U$$929/B sky130_fd_sc_hd__buf_6
XFILLER_107_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1289 U$$3697/B VGND VGND VPWR VPWR U$$3698/A sky130_fd_sc_hd__buf_6
XFILLER_4_395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4469_1811 VGND VGND VPWR VPWR U$$4469_1811/HI U$$4469/B sky130_fd_sc_hd__conb_1
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_328 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$890 U$$890/A1 U$$892/A2 U$$892/A1 U$$892/B2 VGND VGND VPWR VPWR U$$891/A sky130_fd_sc_hd__a22o_1
XFILLER_91_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1040 U$$1040/A U$$980/B VGND VGND VPWR VPWR U$$1040/X sky130_fd_sc_hd__xor2_1
XU$$1051 U$$914/A1 U$$965/A2 U$$914/B1 U$$965/B2 VGND VGND VPWR VPWR U$$1052/A sky130_fd_sc_hd__a22o_1
XFILLER_91_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1062 U$$1062/A U$$994/B VGND VGND VPWR VPWR U$$1062/X sky130_fd_sc_hd__xor2_1
XFILLER_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1073 U$$799/A1 U$$1093/A2 U$$938/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1074/A sky130_fd_sc_hd__a22o_1
XFILLER_52_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1084 U$$1084/A U$$1084/B VGND VGND VPWR VPWR U$$1084/X sky130_fd_sc_hd__xor2_1
XFILLER_149_636 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1095 U$$1095/A VGND VGND VPWR VPWR U$$1095/Y sky130_fd_sc_hd__inv_1
XFILLER_177_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1076 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_81_6 U$$3627/X U$$3760/X U$$3893/X VGND VGND VPWR VPWR dadda_fa_2_82_3/A
+ dadda_fa_2_81_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_74_5 U$$3746/X U$$3879/X U$$4012/X VGND VGND VPWR VPWR dadda_fa_2_75_2/A
+ dadda_fa_2_74_5/A sky130_fd_sc_hd__fa_1
XFILLER_86_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_67_4 U$$4131/X U$$4264/X U$$4397/X VGND VGND VPWR VPWR dadda_fa_2_68_1/CIN
+ dadda_fa_2_67_4/CIN sky130_fd_sc_hd__fa_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_37_2 dadda_fa_4_37_2/A dadda_fa_4_37_2/B dadda_fa_4_37_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_38_0/CIN dadda_fa_5_37_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_54_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_25 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_831 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_63_5 U$$2128/X U$$2261/X VGND VGND VPWR VPWR dadda_fa_1_64_7/A dadda_fa_2_63_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_118_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_62_3 U$$1328/X U$$1461/X U$$1594/X VGND VGND VPWR VPWR dadda_fa_1_63_6/B
+ dadda_fa_1_62_8/B sky130_fd_sc_hd__fa_1
XTAP_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3904 U$$4176/B1 U$$3840/X U$$4043/A1 U$$3841/X VGND VGND VPWR VPWR U$$3905/A sky130_fd_sc_hd__a22o_1
XU$$3915 U$$3915/A U$$3967/B VGND VGND VPWR VPWR U$$3915/X sky130_fd_sc_hd__xor2_1
XU$$3926 U$$912/A1 U$$3926/A2 U$$4476/A1 U$$3926/B2 VGND VGND VPWR VPWR U$$3927/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3937 U$$3937/A U$$3967/B VGND VGND VPWR VPWR U$$3937/X sky130_fd_sc_hd__xor2_1
XTAP_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$270 final_adder.U$$272/B final_adder.U$$270/B VGND VGND VPWR VPWR
+ final_adder.U$$396/B sky130_fd_sc_hd__and2_1
XTAP_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3948 U$$521/B1 U$$3966/A2 U$$4498/A1 U$$3966/B2 VGND VGND VPWR VPWR U$$3949/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$281 final_adder.U$$280/B final_adder.U$$155/X final_adder.U$$153/X
+ VGND VGND VPWR VPWR final_adder.U$$281/X sky130_fd_sc_hd__a21o_1
XTAP_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_32_1 dadda_fa_3_32_1/A dadda_fa_3_32_1/B dadda_fa_3_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_0/CIN dadda_fa_4_32_2/A sky130_fd_sc_hd__fa_1
XU$$120 U$$942/A1 U$$122/A2 U$$122/A1 U$$122/B2 VGND VGND VPWR VPWR U$$121/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$292 final_adder.U$$294/B final_adder.U$$292/B VGND VGND VPWR VPWR
+ final_adder.U$$418/B sky130_fd_sc_hd__and2_1
XU$$3959 U$$3959/A U$$3972/A VGND VGND VPWR VPWR U$$3959/X sky130_fd_sc_hd__xor2_1
XTAP_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$131 U$$131/A U$$99/B VGND VGND VPWR VPWR U$$131/X sky130_fd_sc_hd__xor2_1
XFILLER_166_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$142 U$$140/B U$$136/A U$$138/A U$$137/Y VGND VGND VPWR VPWR U$$142/X sky130_fd_sc_hd__a22o_4
XTAP_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$153 U$$16/A1 U$$175/A2 U$$18/A1 U$$175/B2 VGND VGND VPWR VPWR U$$154/A sky130_fd_sc_hd__a22o_1
XTAP_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$164 U$$164/A U$$184/B VGND VGND VPWR VPWR U$$164/X sky130_fd_sc_hd__xor2_1
XTAP_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_25_0 U$$722/X U$$855/X U$$988/X VGND VGND VPWR VPWR dadda_fa_4_26_0/B
+ dadda_fa_4_25_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$175 U$$38/A1 U$$175/A2 U$$40/A1 U$$175/B2 VGND VGND VPWR VPWR U$$176/A sky130_fd_sc_hd__a22o_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$186 U$$186/A U$$212/B VGND VGND VPWR VPWR U$$186/X sky130_fd_sc_hd__xor2_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$197 U$$882/A1 U$$217/A2 U$$882/B1 U$$217/B2 VGND VGND VPWR VPWR U$$198/A sky130_fd_sc_hd__a22o_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4499_1826 VGND VGND VPWR VPWR U$$4499_1826/HI U$$4499/B sky130_fd_sc_hd__conb_1
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_398_ _399_/CLK _398_/D VGND VGND VPWR VPWR _398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_91_5 dadda_fa_2_91_5/A dadda_fa_2_91_5/B dadda_fa_2_91_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_92_2/A dadda_fa_4_91_0/A sky130_fd_sc_hd__fa_2
Xrepeater1020 input86/X VGND VGND VPWR VPWR U$$3078/B1 sky130_fd_sc_hd__buf_6
Xrepeater1031 input85/X VGND VGND VPWR VPWR U$$4311/A1 sky130_fd_sc_hd__buf_6
XFILLER_86_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1042 U$$2661/B1 VGND VGND VPWR VPWR U$$60/A1 sky130_fd_sc_hd__buf_4
XFILLER_99_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1053 U$$3207/B1 VGND VGND VPWR VPWR U$$56/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_84_4 dadda_fa_2_84_4/A dadda_fa_2_84_4/B dadda_fa_2_84_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_1/CIN dadda_fa_3_84_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1064 input81/X VGND VGND VPWR VPWR U$$4029/A1 sky130_fd_sc_hd__buf_6
XFILLER_142_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1075 U$$3612/B1 VGND VGND VPWR VPWR U$$52/A1 sky130_fd_sc_hd__buf_4
Xrepeater1086 U$$3884/B1 VGND VGND VPWR VPWR U$$2925/B1 sky130_fd_sc_hd__buf_4
XFILLER_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1097 input77/X VGND VGND VPWR VPWR U$$4293/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_77_3 dadda_fa_2_77_3/A dadda_fa_2_77_3/B dadda_fa_2_77_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/B dadda_fa_3_77_3/B sky130_fd_sc_hd__fa_1
XFILLER_141_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_47_1 dadda_fa_5_47_1/A dadda_fa_5_47_1/B dadda_fa_5_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_48_0/B dadda_fa_7_47_0/A sky130_fd_sc_hd__fa_1
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_100_2 U$$3266/X U$$3399/X U$$3532/X VGND VGND VPWR VPWR dadda_fa_3_101_2/A
+ dadda_fa_3_100_3/B sky130_fd_sc_hd__fa_1
XFILLER_63_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_121_1 dadda_fa_5_121_1/A dadda_fa_5_121_1/B dadda_fa_5_121_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_122_0/B dadda_fa_7_121_0/A sky130_fd_sc_hd__fa_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_114_0 dadda_fa_5_114_0/A dadda_fa_5_114_0/B dadda_fa_5_114_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_115_0/A dadda_fa_6_114_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_191_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_992 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_72_2 U$$2811/X U$$2944/X U$$3077/X VGND VGND VPWR VPWR dadda_fa_2_73_1/A
+ dadda_fa_2_72_4/A sky130_fd_sc_hd__fa_1
XFILLER_120_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_65_1 U$$2930/X U$$3063/X U$$3196/X VGND VGND VPWR VPWR dadda_fa_2_66_0/CIN
+ dadda_fa_2_65_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_42_0 dadda_fa_4_42_0/A dadda_fa_4_42_0/B dadda_fa_4_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/A dadda_fa_5_42_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_58_0 U$$1586/X U$$1719/X U$$1852/X VGND VGND VPWR VPWR dadda_fa_2_59_0/B
+ dadda_fa_2_58_3/B sky130_fd_sc_hd__fa_1
XFILLER_101_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1809 U$$4410/B1 U$$1831/A2 U$$989/A1 U$$1831/B2 VGND VGND VPWR VPWR U$$1810/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_321_ _329_/CLK _321_/D VGND VGND VPWR VPWR _321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_252_ _255_/CLK _252_/D VGND VGND VPWR VPWR _252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_252 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_183_ _337_/CLK _183_/D VGND VGND VPWR VPWR _183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_94_3 dadda_fa_3_94_3/A dadda_fa_3_94_3/B dadda_fa_3_94_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_95_1/B dadda_fa_4_94_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_202_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_87_2 dadda_fa_3_87_2/A dadda_fa_3_87_2/B dadda_fa_3_87_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_1/A dadda_fa_4_87_2/B sky130_fd_sc_hd__fa_1
XFILLER_135_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_0_54_1 U$$514/X U$$647/X VGND VGND VPWR VPWR dadda_fa_1_55_8/B dadda_fa_2_54_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_123_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_57_0 dadda_fa_6_57_0/A dadda_fa_6_57_0/B dadda_fa_6_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_58_0/B dadda_fa_7_57_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_81_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater709 U$$3841/X VGND VGND VPWR VPWR U$$3968/B2 sky130_fd_sc_hd__buf_8
XU$$4402 U$$4402/A1 U$$4388/X U$$4402/B1 U$$4432/B2 VGND VGND VPWR VPWR U$$4403/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4413 U$$4413/A U$$4413/B VGND VGND VPWR VPWR U$$4413/X sky130_fd_sc_hd__xor2_1
XFILLER_38_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_60_0 U$$127/X U$$260/X U$$393/X VGND VGND VPWR VPWR dadda_fa_1_61_6/A
+ dadda_fa_1_60_7/CIN sky130_fd_sc_hd__fa_1
XU$$4424 U$$4424/A1 U$$4388/X input73/X U$$4426/B2 VGND VGND VPWR VPWR U$$4425/A sky130_fd_sc_hd__a22o_1
XU$$4435 U$$4435/A U$$4435/B VGND VGND VPWR VPWR U$$4435/X sky130_fd_sc_hd__xor2_1
XU$$4446 input84/X U$$4388/X input85/X U$$4498/B2 VGND VGND VPWR VPWR U$$4447/A sky130_fd_sc_hd__a22o_1
XU$$3701 U$$3836/A VGND VGND VPWR VPWR U$$3701/Y sky130_fd_sc_hd__inv_1
XFILLER_92_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3712 U$$3712/A U$$3754/B VGND VGND VPWR VPWR U$$3712/X sky130_fd_sc_hd__xor2_1
XTAP_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_116_2 input147/X dadda_fa_4_116_2/B dadda_ha_3_116_0/SUM VGND VGND VPWR
+ VPWR dadda_fa_5_117_0/CIN dadda_fa_5_116_1/CIN sky130_fd_sc_hd__fa_1
XU$$4457 U$$4457/A U$$4457/B VGND VGND VPWR VPWR U$$4457/X sky130_fd_sc_hd__xor2_1
XU$$4468 input96/X U$$4388/X U$$4468/B1 U$$4486/B2 VGND VGND VPWR VPWR U$$4469/A sky130_fd_sc_hd__a22o_1
XTAP_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3723 U$$4269/B1 U$$3739/A2 U$$4408/B1 U$$3739/B2 VGND VGND VPWR VPWR U$$3724/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4479 U$$4479/A U$$4479/B VGND VGND VPWR VPWR U$$4479/X sky130_fd_sc_hd__xor2_1
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3734 U$$3734/A U$$3740/B VGND VGND VPWR VPWR U$$3734/X sky130_fd_sc_hd__xor2_1
XTAP_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3745 U$$3880/B1 U$$3753/A2 U$$3747/A1 U$$3753/B2 VGND VGND VPWR VPWR U$$3746/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3756 U$$3756/A U$$3778/B VGND VGND VPWR VPWR U$$3756/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_109_1 dadda_fa_4_109_1/A dadda_fa_4_109_1/B dadda_fa_4_109_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/B dadda_fa_5_109_1/B sky130_fd_sc_hd__fa_1
XTAP_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3767 U$$3902/B1 U$$3773/A2 U$$4043/A1 U$$3773/B2 VGND VGND VPWR VPWR U$$3768/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3778 U$$3778/A U$$3778/B VGND VGND VPWR VPWR U$$3778/X sky130_fd_sc_hd__xor2_1
XU$$3789 U$$912/A1 U$$3793/A2 U$$4476/A1 U$$3793/B2 VGND VGND VPWR VPWR U$$3790/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_82_1 dadda_fa_2_82_1/A dadda_fa_2_82_1/B dadda_fa_2_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_0/CIN dadda_fa_3_82_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_75_0 dadda_fa_2_75_0/A dadda_fa_2_75_0/B dadda_fa_2_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_0/B dadda_fa_3_75_2/B sky130_fd_sc_hd__fa_1
XFILLER_130_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_51_7 U$$2902/X U$$3035/X U$$3168/X VGND VGND VPWR VPWR dadda_fa_2_52_2/CIN
+ dadda_fa_2_51_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_97_1 dadda_fa_4_97_1/A dadda_fa_4_97_1/B dadda_fa_4_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/B dadda_fa_5_97_1/B sky130_fd_sc_hd__fa_1
XFILLER_137_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_74_0 dadda_fa_7_74_0/A dadda_fa_7_74_0/B dadda_fa_7_74_0/CIN VGND VGND
+ VPWR VPWR _371_/D _242_/D sky130_fd_sc_hd__fa_2
XFILLER_180_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3008 U$$3008/A U$$3008/B VGND VGND VPWR VPWR U$$3008/X sky130_fd_sc_hd__xor2_1
XFILLER_46_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3019 U$$3017/B input38/X input39/X U$$3014/Y VGND VGND VPWR VPWR U$$3019/X sky130_fd_sc_hd__a22o_2
XFILLER_207_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2307 U$$2307/A U$$2311/B VGND VGND VPWR VPWR U$$2307/X sky130_fd_sc_hd__xor2_1
XFILLER_34_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2318 U$$3960/B1 U$$2326/A2 U$$2318/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2319/A
+ sky130_fd_sc_hd__a22o_1
XU$$2329 input27/X VGND VGND VPWR VPWR U$$2329/Y sky130_fd_sc_hd__inv_1
XFILLER_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1606 U$$1606/A U$$1608/B VGND VGND VPWR VPWR U$$1606/X sky130_fd_sc_hd__xor2_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1617 U$$2165/A1 U$$1635/A2 U$$660/A1 U$$1635/B2 VGND VGND VPWR VPWR U$$1618/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1628 U$$1628/A U$$1628/B VGND VGND VPWR VPWR U$$1628/X sky130_fd_sc_hd__xor2_1
XFILLER_163_1204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1639 U$$4516/A1 U$$1511/X U$$4516/B1 U$$1512/X VGND VGND VPWR VPWR U$$1640/A sky130_fd_sc_hd__a22o_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_304_ _304_/CLK _304_/D VGND VGND VPWR VPWR _304_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_235_ _367_/CLK _235_/D VGND VGND VPWR VPWR _235_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_204_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1002 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_92_0 dadda_fa_3_92_0/A dadda_fa_3_92_0/B dadda_fa_3_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_0/B dadda_fa_4_92_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_13_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater506 U$$3132/A2 VGND VGND VPWR VPWR U$$3124/A2 sky130_fd_sc_hd__buf_6
XFILLER_46_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater517 U$$2881/X VGND VGND VPWR VPWR U$$2977/A2 sky130_fd_sc_hd__buf_4
XFILLER_78_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4210 U$$4210/A1 U$$4210/A2 U$$4210/B1 U$$4210/B2 VGND VGND VPWR VPWR U$$4211/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater528 U$$2810/A2 VGND VGND VPWR VPWR U$$2796/A2 sky130_fd_sc_hd__buf_4
XFILLER_78_784 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4221 U$$4221/A U$$4247/A VGND VGND VPWR VPWR U$$4221/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_54_5 dadda_fa_2_54_5/A dadda_fa_2_54_5/B dadda_fa_2_54_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_55_2/A dadda_fa_4_54_0/A sky130_fd_sc_hd__fa_1
XFILLER_133_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater539 U$$2711/A2 VGND VGND VPWR VPWR U$$2691/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_121_0 U$$3972/Y U$$4106/X U$$4239/X VGND VGND VPWR VPWR dadda_fa_5_122_1/B
+ dadda_fa_5_121_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4232 U$$4506/A1 U$$4238/A2 U$$4369/B1 U$$4238/B2 VGND VGND VPWR VPWR U$$4233/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4243 U$$4243/A U$$4243/B VGND VGND VPWR VPWR U$$4243/X sky130_fd_sc_hd__xor2_1
XU$$4254 U$$4254/A U$$4278/B VGND VGND VPWR VPWR U$$4254/X sky130_fd_sc_hd__xor2_1
XFILLER_65_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3520 U$$3520/A U$$3550/B VGND VGND VPWR VPWR U$$3520/X sky130_fd_sc_hd__xor2_1
XU$$4265 U$$4402/A1 U$$4297/A2 U$$4402/B1 U$$4297/B2 VGND VGND VPWR VPWR U$$4266/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_47_4 dadda_fa_2_47_4/A dadda_fa_2_47_4/B dadda_fa_2_47_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_1/CIN dadda_fa_3_47_3/CIN sky130_fd_sc_hd__fa_1
XU$$3531 U$$4077/B1 U$$3549/A2 U$$3944/A1 U$$3549/B2 VGND VGND VPWR VPWR U$$3532/A
+ sky130_fd_sc_hd__a22o_1
XU$$4276 U$$4276/A U$$4278/B VGND VGND VPWR VPWR U$$4276/X sky130_fd_sc_hd__xor2_1
XFILLER_93_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3542 U$$3542/A U$$3561/A VGND VGND VPWR VPWR U$$3542/X sky130_fd_sc_hd__xor2_1
XFILLER_92_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4287 U$$4424/A1 U$$4297/A2 U$$4289/A1 U$$4297/B2 VGND VGND VPWR VPWR U$$4288/A
+ sky130_fd_sc_hd__a22o_1
XU$$3553 input121/X U$$3559/A2 input122/X U$$3559/B2 VGND VGND VPWR VPWR U$$3554/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4298 U$$4298/A U$$4310/B VGND VGND VPWR VPWR U$$4298/X sky130_fd_sc_hd__xor2_1
XFILLER_81_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3564 U$$3643/B VGND VGND VPWR VPWR U$$3564/Y sky130_fd_sc_hd__inv_1
XU$$3575 U$$3575/A U$$3665/B VGND VGND VPWR VPWR U$$3575/X sky130_fd_sc_hd__xor2_1
XFILLER_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2830 U$$3378/A1 U$$2844/A2 U$$3243/A1 U$$2844/B2 VGND VGND VPWR VPWR U$$2831/A
+ sky130_fd_sc_hd__a22o_1
XU$$2841 U$$2841/A U$$2845/B VGND VGND VPWR VPWR U$$2841/X sky130_fd_sc_hd__xor2_1
XU$$3586 U$$4269/B1 U$$3606/A2 U$$4408/B1 U$$3606/B2 VGND VGND VPWR VPWR U$$3587/A
+ sky130_fd_sc_hd__a22o_1
XU$$2852 U$$521/B1 U$$2858/A2 U$$660/B1 U$$2858/B2 VGND VGND VPWR VPWR U$$2853/A sky130_fd_sc_hd__a22o_1
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3597 U$$3597/A U$$3637/B VGND VGND VPWR VPWR U$$3597/X sky130_fd_sc_hd__xor2_1
XU$$2863 U$$2863/A U$$2869/B VGND VGND VPWR VPWR U$$2863/X sky130_fd_sc_hd__xor2_1
XU$$2874 U$$3557/B1 U$$2874/A2 U$$2874/B1 U$$2874/B2 VGND VGND VPWR VPWR U$$2875/A
+ sky130_fd_sc_hd__a22o_1
XU$$2885 U$$3159/A1 U$$2921/A2 U$$3159/B1 U$$2921/B2 VGND VGND VPWR VPWR U$$2886/A
+ sky130_fd_sc_hd__a22o_1
XU$$2896 U$$2896/A U$$2922/B VGND VGND VPWR VPWR U$$2896/X sky130_fd_sc_hd__xor2_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_190 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_209_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$803 final_adder.U$$770/A final_adder.U$$723/X final_adder.U$$691/X
+ VGND VGND VPWR VPWR final_adder.U$$803/X sky130_fd_sc_hd__a21o_1
XFILLER_190_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$825 final_adder.U$$792/A final_adder.U$$625/X final_adder.U$$713/X
+ VGND VGND VPWR VPWR final_adder.U$$825/X sky130_fd_sc_hd__a21o_1
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$847 final_adder.U$$750/X final_adder.U$$815/X final_adder.U$$751/X
+ VGND VGND VPWR VPWR final_adder.U$$847/X sky130_fd_sc_hd__a21o_2
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$869 final_adder.U$$772/X final_adder.U$$725/X final_adder.U$$773/X
+ VGND VGND VPWR VPWR final_adder.U$$869/X sky130_fd_sc_hd__a21o_2
XU$$708 U$$708/A U$$740/B VGND VGND VPWR VPWR U$$708/X sky130_fd_sc_hd__xor2_1
XFILLER_72_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$719 U$$854/B1 U$$739/A2 U$$719/B1 U$$739/B2 VGND VGND VPWR VPWR U$$720/A sky130_fd_sc_hd__a22o_1
XFILLER_16_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_42_3 U$$1288/X U$$1421/X U$$1554/X VGND VGND VPWR VPWR dadda_fa_2_43_4/A
+ dadda_fa_2_42_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_186_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_12_1 U$$430/X U$$563/X U$$696/X VGND VGND VPWR VPWR dadda_fa_5_13_0/B
+ dadda_fa_5_12_1/B sky130_fd_sc_hd__fa_1
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_634 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$143_1717 VGND VGND VPWR VPWR U$$143_1717/HI U$$143/A1 sky130_fd_sc_hd__conb_1
XFILLER_71_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1608 U$$4494/A1 VGND VGND VPWR VPWR U$$2165/A1 sky130_fd_sc_hd__buf_4
XFILLER_180_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1619 U$$1370/A VGND VGND VPWR VPWR U$$1354/B sky130_fd_sc_hd__buf_8
XFILLER_153_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_109_0 U$$3150/Y U$$3284/X U$$3417/X VGND VGND VPWR VPWR dadda_fa_4_110_0/B
+ dadda_fa_4_109_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_57_3 dadda_fa_3_57_3/A dadda_fa_3_57_3/B dadda_fa_3_57_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_58_1/B dadda_fa_4_57_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2104 U$$2104/A U$$2114/B VGND VGND VPWR VPWR U$$2104/X sky130_fd_sc_hd__xor2_1
XFILLER_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2115 U$$3483/B1 U$$2189/A2 input84/X U$$2189/B2 VGND VGND VPWR VPWR U$$2116/A
+ sky130_fd_sc_hd__a22o_1
XU$$2126 U$$2126/A U$$2170/B VGND VGND VPWR VPWR U$$2126/X sky130_fd_sc_hd__xor2_1
XU$$2137 U$$3368/B1 U$$2169/A2 U$$3235/A1 U$$2169/B2 VGND VGND VPWR VPWR U$$2138/A
+ sky130_fd_sc_hd__a22o_1
XU$$2148 U$$2148/A U$$2184/B VGND VGND VPWR VPWR U$$2148/X sky130_fd_sc_hd__xor2_1
XU$$1403 U$$1403/A U$$1405/B VGND VGND VPWR VPWR U$$1403/X sky130_fd_sc_hd__xor2_1
XU$$1414 U$$864/B1 U$$1422/A2 U$$594/A1 U$$1422/B2 VGND VGND VPWR VPWR U$$1415/A sky130_fd_sc_hd__a22o_1
XU$$2159 U$$2568/B1 U$$2183/A2 U$$2159/B1 U$$2183/B2 VGND VGND VPWR VPWR U$$2160/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_612 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1425 U$$1425/A U$$1459/B VGND VGND VPWR VPWR U$$1425/X sky130_fd_sc_hd__xor2_1
XFILLER_76_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1436 U$$1984/A1 U$$1448/A2 U$$342/A1 U$$1448/B2 VGND VGND VPWR VPWR U$$1437/A
+ sky130_fd_sc_hd__a22o_1
XU$$1447 U$$1447/A U$$1449/B VGND VGND VPWR VPWR U$$1447/X sky130_fd_sc_hd__xor2_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1458 U$$2415/B1 U$$1462/A2 U$$90/A1 U$$1462/B2 VGND VGND VPWR VPWR U$$1459/A sky130_fd_sc_hd__a22o_1
XFILLER_203_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1469 U$$1469/A U$$1506/A VGND VGND VPWR VPWR U$$1469/X sky130_fd_sc_hd__xor2_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_218_ _218_/CLK _218_/D VGND VGND VPWR VPWR _218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_450 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4253_1764 VGND VGND VPWR VPWR U$$4253_1764/HI U$$4253/A1 sky130_fd_sc_hd__conb_1
XFILLER_211_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_52_2 dadda_fa_2_52_2/A dadda_fa_2_52_2/B dadda_fa_2_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/A dadda_fa_3_52_3/A sky130_fd_sc_hd__fa_1
XFILLER_66_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4040 U$$4040/A U$$4109/A VGND VGND VPWR VPWR U$$4040/X sky130_fd_sc_hd__xor2_1
XFILLER_211_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4051 input93/X U$$4079/A2 U$$4464/A1 U$$4079/B2 VGND VGND VPWR VPWR U$$4052/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_45_1 U$$2757/X U$$2890/X U$$3023/X VGND VGND VPWR VPWR dadda_fa_3_46_0/CIN
+ dadda_fa_3_45_2/CIN sky130_fd_sc_hd__fa_1
XU$$4062 U$$4062/A U$$4078/B VGND VGND VPWR VPWR U$$4062/X sky130_fd_sc_hd__xor2_1
XU$$4073 U$$4210/A1 U$$4077/A2 U$$4210/B1 U$$4077/B2 VGND VGND VPWR VPWR U$$4074/A
+ sky130_fd_sc_hd__a22o_1
XU$$4084 U$$4084/A U$$4110/A VGND VGND VPWR VPWR U$$4084/X sky130_fd_sc_hd__xor2_1
XU$$4095 U$$4095/A1 U$$4103/A2 U$$4369/B1 U$$4103/B2 VGND VGND VPWR VPWR U$$4096/A
+ sky130_fd_sc_hd__a22o_1
XU$$3350 input84/X U$$3394/A2 input85/X U$$3390/B2 VGND VGND VPWR VPWR U$$3351/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_22_0 dadda_fa_5_22_0/A dadda_fa_5_22_0/B dadda_fa_5_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_23_0/A dadda_fa_6_22_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_38_0 U$$1147/X U$$1280/X U$$1413/X VGND VGND VPWR VPWR dadda_fa_3_39_0/B
+ dadda_fa_3_38_2/B sky130_fd_sc_hd__fa_1
XU$$3361 U$$3361/A U$$3425/A VGND VGND VPWR VPWR U$$3361/X sky130_fd_sc_hd__xor2_1
XFILLER_207_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3372 U$$3644/B1 U$$3374/A2 U$$3511/A1 U$$3374/B2 VGND VGND VPWR VPWR U$$3373/A
+ sky130_fd_sc_hd__a22o_1
XU$$3383 U$$3383/A U$$3417/B VGND VGND VPWR VPWR U$$3383/X sky130_fd_sc_hd__xor2_1
XU$$3394 U$$4077/B1 U$$3394/A2 U$$3944/A1 U$$3394/B2 VGND VGND VPWR VPWR U$$3395/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2660 U$$2660/A U$$2680/B VGND VGND VPWR VPWR U$$2660/X sky130_fd_sc_hd__xor2_1
XU$$2671 U$$3902/B1 U$$2711/A2 U$$2808/B1 U$$2711/B2 VGND VGND VPWR VPWR U$$2672/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2682 U$$2682/A U$$2716/B VGND VGND VPWR VPWR U$$2682/X sky130_fd_sc_hd__xor2_1
XFILLER_61_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2693 U$$3378/A1 U$$2737/A2 U$$3517/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2694/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1970 U$$3749/B1 U$$1970/A2 U$$52/B1 U$$1970/B2 VGND VGND VPWR VPWR U$$1971/A sky130_fd_sc_hd__a22o_1
XU$$1981 U$$1981/A U$$2017/B VGND VGND VPWR VPWR U$$1981/X sky130_fd_sc_hd__xor2_1
XFILLER_166_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1992 U$$896/A1 U$$2040/A2 U$$759/B1 U$$2040/B2 VGND VGND VPWR VPWR U$$1993/A sky130_fd_sc_hd__a22o_1
XFILLER_142_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_67_2 dadda_fa_4_67_2/A dadda_fa_4_67_2/B dadda_fa_4_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_68_0/CIN dadda_fa_5_67_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput106 b[47] VGND VGND VPWR VPWR input106/X sky130_fd_sc_hd__buf_6
Xinput117 b[57] VGND VGND VPWR VPWR input117/X sky130_fd_sc_hd__buf_6
Xinput128 b[9] VGND VGND VPWR VPWR input128/X sky130_fd_sc_hd__buf_6
XTAP_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput139 c[109] VGND VGND VPWR VPWR input139/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$600 final_adder.U$$608/B final_adder.U$$600/B VGND VGND VPWR VPWR
+ final_adder.U$$720/B sky130_fd_sc_hd__and2_1
XTAP_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$611 final_adder.U$$610/B final_adder.U$$495/X final_adder.U$$487/X
+ VGND VGND VPWR VPWR final_adder.U$$611/X sky130_fd_sc_hd__a21o_1
XTAP_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_37_0 dadda_fa_7_37_0/A dadda_fa_7_37_0/B dadda_fa_7_37_0/CIN VGND VGND
+ VPWR VPWR _334_/D _205_/D sky130_fd_sc_hd__fa_2
XFILLER_5_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$633 final_adder.U$$632/B final_adder.U$$529/X final_adder.U$$513/X
+ VGND VGND VPWR VPWR final_adder.U$$633/X sky130_fd_sc_hd__a21o_1
XTAP_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$644 final_adder.U$$660/B final_adder.U$$644/B VGND VGND VPWR VPWR
+ final_adder.U$$756/B sky130_fd_sc_hd__and2_1
XTAP_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$655 final_adder.U$$654/B final_adder.U$$551/X final_adder.U$$535/X
+ VGND VGND VPWR VPWR final_adder.U$$655/X sky130_fd_sc_hd__a21o_1
XTAP_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$666 final_adder.U$$682/B final_adder.U$$666/B VGND VGND VPWR VPWR
+ final_adder.U$$778/B sky130_fd_sc_hd__and2_1
XTAP_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater870 U$$1375/X VGND VGND VPWR VPWR U$$1504/B2 sky130_fd_sc_hd__buf_8
XU$$505 U$$916/A1 U$$521/A2 U$$916/B1 U$$521/B2 VGND VGND VPWR VPWR U$$506/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$677 final_adder.U$$676/B final_adder.U$$573/X final_adder.U$$557/X
+ VGND VGND VPWR VPWR final_adder.U$$677/X sky130_fd_sc_hd__a21o_1
XFILLER_186_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$516 U$$516/A U$$516/B VGND VGND VPWR VPWR U$$516/X sky130_fd_sc_hd__xor2_1
XFILLER_5_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_40_0 U$$87/X U$$220/X U$$353/X VGND VGND VPWR VPWR dadda_fa_2_41_3/CIN
+ dadda_fa_2_40_5/A sky130_fd_sc_hd__fa_1
Xrepeater881 U$$1190/B2 VGND VGND VPWR VPWR U$$1174/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$688 final_adder.U$$704/B final_adder.U$$688/B VGND VGND VPWR VPWR
+ final_adder.U$$800/B sky130_fd_sc_hd__and2_1
XTAP_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$527 U$$527/A1 U$$527/A2 U$$527/B1 U$$527/B2 VGND VGND VPWR VPWR U$$528/A sky130_fd_sc_hd__a22o_1
XFILLER_56_275 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater892 U$$134/B2 VGND VGND VPWR VPWR U$$122/B2 sky130_fd_sc_hd__buf_8
Xfinal_adder.U$$699 final_adder.U$$698/B final_adder.U$$595/X final_adder.U$$579/X
+ VGND VGND VPWR VPWR final_adder.U$$699/X sky130_fd_sc_hd__a21o_1
XU$$538 U$$538/A U$$546/B VGND VGND VPWR VPWR U$$538/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$549 U$$549/A VGND VGND VPWR VPWR U$$551/B sky130_fd_sc_hd__inv_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1405 U$$2170/B VGND VGND VPWR VPWR U$$2092/B sky130_fd_sc_hd__buf_6
XFILLER_126_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1416 U$$2037/B VGND VGND VPWR VPWR U$$2009/B sky130_fd_sc_hd__buf_8
XFILLER_125_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1427 input20/X VGND VGND VPWR VPWR U$$1914/B sky130_fd_sc_hd__buf_6
XFILLER_125_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1438 U$$1620/B VGND VGND VPWR VPWR U$$1574/B sky130_fd_sc_hd__buf_6
XFILLER_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1449 U$$1506/A VGND VGND VPWR VPWR U$$1459/B sky130_fd_sc_hd__buf_8
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_62_1 dadda_fa_3_62_1/A dadda_fa_3_62_1/B dadda_fa_3_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_0/CIN dadda_fa_4_62_2/A sky130_fd_sc_hd__fa_1
XFILLER_0_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_55_0 dadda_fa_3_55_0/A dadda_fa_3_55_0/B dadda_fa_3_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_0/B dadda_fa_4_55_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1200 U$$2842/B1 U$$1204/A2 U$$2709/A1 U$$1204/B2 VGND VGND VPWR VPWR U$$1201/A
+ sky130_fd_sc_hd__a22o_1
XU$$1211 U$$1211/A U$$1232/A VGND VGND VPWR VPWR U$$1211/X sky130_fd_sc_hd__xor2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1222 U$$3414/A1 U$$1222/A2 U$$3414/B1 U$$1222/B2 VGND VGND VPWR VPWR U$$1223/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1233 input9/X VGND VGND VPWR VPWR U$$1233/Y sky130_fd_sc_hd__inv_1
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1244 U$$1244/A U$$1272/B VGND VGND VPWR VPWR U$$1244/X sky130_fd_sc_hd__xor2_1
XU$$1255 U$$1666/A1 U$$1289/A2 U$$1666/B1 U$$1281/B2 VGND VGND VPWR VPWR U$$1256/A
+ sky130_fd_sc_hd__a22o_1
XU$$1266 U$$1266/A U$$1270/B VGND VGND VPWR VPWR U$$1266/X sky130_fd_sc_hd__xor2_1
XU$$1277 U$$864/B1 U$$1323/A2 U$$731/A1 U$$1307/B2 VGND VGND VPWR VPWR U$$1278/A sky130_fd_sc_hd__a22o_1
XU$$1288 U$$1288/A U$$1330/B VGND VGND VPWR VPWR U$$1288/X sky130_fd_sc_hd__xor2_1
XU$$1299 U$$477/A1 U$$1323/A2 U$$342/A1 U$$1307/B2 VGND VGND VPWR VPWR U$$1300/A sky130_fd_sc_hd__a22o_1
XFILLER_30_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_112_0 dadda_fa_7_112_0/A dadda_fa_7_112_0/B dadda_fa_7_112_0/CIN VGND
+ VGND VPWR VPWR _409_/D _280_/D sky130_fd_sc_hd__fa_1
XFILLER_129_531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1060 final_adder.U$$218/A final_adder.U$$831/X VGND VGND VPWR VPWR
+ output314/A sky130_fd_sc_hd__xor2_1
XFILLER_144_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1071 final_adder.U$$208/B final_adder.U$$979/X VGND VGND VPWR VPWR
+ output326/A sky130_fd_sc_hd__xor2_1
XFILLER_7_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1082 final_adder.U$$196/A final_adder.U$$809/X VGND VGND VPWR VPWR
+ output338/A sky130_fd_sc_hd__xor2_1
XFILLER_144_556 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1093 final_adder.U$$186/B final_adder.U$$957/X VGND VGND VPWR VPWR
+ output350/A sky130_fd_sc_hd__xor2_1
XFILLER_172_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_77_1 dadda_fa_5_77_1/A dadda_fa_5_77_1/B dadda_fa_5_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_78_0/B dadda_fa_7_77_0/A sky130_fd_sc_hd__fa_1
XFILLER_144_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_69_8 dadda_fa_1_69_8/A dadda_fa_1_69_8/B dadda_fa_1_69_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_70_3/A dadda_fa_3_69_0/A sky130_fd_sc_hd__fa_1
XFILLER_97_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4411_1782 VGND VGND VPWR VPWR U$$4411_1782/HI U$$4411/B sky130_fd_sc_hd__conb_1
XFILLER_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3180 U$$3180/A U$$3228/B VGND VGND VPWR VPWR U$$3180/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_9_0 dadda_fa_6_9_0/A dadda_fa_6_9_0/B dadda_fa_6_9_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_10_0/B dadda_fa_7_9_0/CIN sky130_fd_sc_hd__fa_1
XU$$3191 U$$860/B1 U$$3207/A2 U$$3876/B1 U$$3207/B2 VGND VGND VPWR VPWR U$$3192/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2490 U$$2625/B1 U$$2490/A2 U$$2492/A1 U$$2490/B2 VGND VGND VPWR VPWR U$$2491/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_504 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_72_0 dadda_fa_4_72_0/A dadda_fa_4_72_0/B dadda_fa_4_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/A dadda_fa_5_72_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_88_0 dadda_fa_1_88_0/A U$$1779/X U$$1912/X VGND VGND VPWR VPWR dadda_fa_2_89_3/B
+ dadda_fa_2_88_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$430 final_adder.U$$434/B final_adder.U$$430/B VGND VGND VPWR VPWR
+ final_adder.U$$554/B sky130_fd_sc_hd__and2_1
XTAP_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$441 final_adder.U$$440/B final_adder.U$$319/X final_adder.U$$315/X
+ VGND VGND VPWR VPWR final_adder.U$$441/X sky130_fd_sc_hd__a21o_1
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$452 final_adder.U$$456/B final_adder.U$$452/B VGND VGND VPWR VPWR
+ final_adder.U$$576/B sky130_fd_sc_hd__and2_1
XTAP_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$463 final_adder.U$$462/B final_adder.U$$341/X final_adder.U$$337/X
+ VGND VGND VPWR VPWR final_adder.U$$463/X sky130_fd_sc_hd__a21o_1
XTAP_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$302 U$$28/A1 U$$302/A2 U$$578/A1 U$$302/B2 VGND VGND VPWR VPWR U$$303/A sky130_fd_sc_hd__a22o_1
XTAP_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$474 final_adder.U$$478/B final_adder.U$$474/B VGND VGND VPWR VPWR
+ final_adder.U$$598/B sky130_fd_sc_hd__and2_1
XTAP_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$313 U$$313/A U$$343/B VGND VGND VPWR VPWR U$$313/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$485 final_adder.U$$484/B final_adder.U$$363/X final_adder.U$$359/X
+ VGND VGND VPWR VPWR final_adder.U$$485/X sky130_fd_sc_hd__a21o_1
XTAP_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$324 U$$461/A1 U$$350/A2 U$$461/B1 U$$350/B2 VGND VGND VPWR VPWR U$$325/A sky130_fd_sc_hd__a22o_1
XFILLER_84_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$496 final_adder.U$$500/B final_adder.U$$496/B VGND VGND VPWR VPWR
+ final_adder.U$$612/A sky130_fd_sc_hd__and2_1
XTAP_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$335 U$$335/A U$$367/B VGND VGND VPWR VPWR U$$335/X sky130_fd_sc_hd__xor2_1
XFILLER_83_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$346 U$$757/A1 U$$366/A2 U$$483/B1 U$$366/B2 VGND VGND VPWR VPWR U$$347/A sky130_fd_sc_hd__a22o_1
XTAP_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$357 U$$357/A U$$397/B VGND VGND VPWR VPWR U$$357/X sky130_fd_sc_hd__xor2_1
XFILLER_72_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$368 U$$916/A1 U$$378/A2 U$$916/B1 U$$378/B2 VGND VGND VPWR VPWR U$$369/A sky130_fd_sc_hd__a22o_1
XU$$379 U$$379/A U$$379/B VGND VGND VPWR VPWR U$$379/X sky130_fd_sc_hd__xor2_1
XFILLER_16_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_87_0 dadda_fa_6_87_0/A dadda_fa_6_87_0/B dadda_fa_6_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_88_0/B dadda_fa_7_87_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1202 input65/X VGND VGND VPWR VPWR U$$2609/B1 sky130_fd_sc_hd__buf_4
Xrepeater1213 U$$683/B VGND VGND VPWR VPWR U$$685/A sky130_fd_sc_hd__buf_6
Xrepeater1224 U$$4310/B VGND VGND VPWR VPWR U$$4294/B sky130_fd_sc_hd__buf_6
Xrepeater1235 U$$4227/B VGND VGND VPWR VPWR U$$4211/B sky130_fd_sc_hd__clkbuf_8
XFILLER_154_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1246 U$$367/B VGND VGND VPWR VPWR U$$377/B sky130_fd_sc_hd__buf_6
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1257 input55/X VGND VGND VPWR VPWR U$$4110/A sky130_fd_sc_hd__buf_8
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1268 U$$3778/B VGND VGND VPWR VPWR U$$3754/B sky130_fd_sc_hd__buf_8
Xrepeater1279 U$$883/B VGND VGND VPWR VPWR U$$877/B sky130_fd_sc_hd__buf_6
XFILLER_153_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_315 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_811 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$880 U$$56/B1 U$$882/A2 U$$882/A1 U$$882/B2 VGND VGND VPWR VPWR U$$881/A sky130_fd_sc_hd__a22o_1
XU$$1030 U$$1030/A U$$1076/B VGND VGND VPWR VPWR U$$1030/X sky130_fd_sc_hd__xor2_1
XFILLER_17_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$891 U$$891/A U$$929/B VGND VGND VPWR VPWR U$$891/X sky130_fd_sc_hd__xor2_1
XFILLER_211_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1041 U$$82/A1 U$$965/A2 U$$84/A1 U$$965/B2 VGND VGND VPWR VPWR U$$1042/A sky130_fd_sc_hd__a22o_1
XU$$1052 U$$1052/A U$$968/B VGND VGND VPWR VPWR U$$1052/X sky130_fd_sc_hd__xor2_1
XFILLER_189_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1063 U$$926/A1 U$$1083/A2 U$$928/A1 U$$1083/B2 VGND VGND VPWR VPWR U$$1064/A sky130_fd_sc_hd__a22o_1
XFILLER_91_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1074 U$$1074/A U$$1076/B VGND VGND VPWR VPWR U$$1074/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1085 U$$811/A1 U$$1093/A2 U$$2318/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1086/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1096 U$$962/A VGND VGND VPWR VPWR U$$1096/Y sky130_fd_sc_hd__inv_1
XFILLER_149_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4441_1797 VGND VGND VPWR VPWR U$$4441_1797/HI U$$4441/B sky130_fd_sc_hd__conb_1
XFILLER_136_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1030 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4517_1835 VGND VGND VPWR VPWR U$$4517_1835/HI U$$4517/B sky130_fd_sc_hd__conb_1
XFILLER_208_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_81_7 U$$4026/X U$$4159/X U$$4292/X VGND VGND VPWR VPWR dadda_fa_2_82_3/B
+ dadda_fa_3_81_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_74_6 U$$4145/X U$$4278/X U$$4411/X VGND VGND VPWR VPWR dadda_fa_2_75_2/B
+ dadda_fa_2_74_5/B sky130_fd_sc_hd__fa_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_935 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_67_5 input220/X dadda_fa_1_67_5/B dadda_fa_1_67_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_68_2/A dadda_fa_2_67_5/A sky130_fd_sc_hd__fa_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_62_4 U$$1727/X U$$1860/X U$$1993/X VGND VGND VPWR VPWR dadda_fa_1_63_6/CIN
+ dadda_fa_1_62_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3905 U$$3905/A U$$3909/B VGND VGND VPWR VPWR U$$3905/X sky130_fd_sc_hd__xor2_1
XFILLER_44_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3916 U$$4464/A1 U$$3926/A2 U$$4466/A1 U$$3926/B2 VGND VGND VPWR VPWR U$$3917/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_19_2 U$$843/X U$$976/X VGND VGND VPWR VPWR dadda_fa_4_20_1/B dadda_ha_3_19_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_18_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$260 final_adder.U$$262/B final_adder.U$$260/B VGND VGND VPWR VPWR
+ final_adder.U$$386/B sky130_fd_sc_hd__and2_1
XU$$3927 U$$3927/A U$$3927/B VGND VGND VPWR VPWR U$$3927/X sky130_fd_sc_hd__xor2_1
XTAP_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3938 input106/X U$$3968/A2 input107/X U$$3968/B2 VGND VGND VPWR VPWR U$$3939/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$110 U$$521/A1 U$$122/A2 U$$384/B1 U$$122/B2 VGND VGND VPWR VPWR U$$111/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$271 final_adder.U$$270/B final_adder.U$$145/X final_adder.U$$143/X
+ VGND VGND VPWR VPWR final_adder.U$$271/X sky130_fd_sc_hd__a21o_1
XFILLER_206_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3949 U$$3949/A U$$3967/B VGND VGND VPWR VPWR U$$3949/X sky130_fd_sc_hd__xor2_1
XTAP_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$282 final_adder.U$$284/B final_adder.U$$282/B VGND VGND VPWR VPWR
+ final_adder.U$$408/B sky130_fd_sc_hd__and2_1
XTAP_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_32_2 dadda_fa_3_32_2/A dadda_fa_3_32_2/B dadda_fa_3_32_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_1/A dadda_fa_4_32_2/B sky130_fd_sc_hd__fa_1
XU$$121 U$$121/A U$$127/B VGND VGND VPWR VPWR U$$121/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$293 final_adder.U$$292/B final_adder.U$$167/X final_adder.U$$165/X
+ VGND VGND VPWR VPWR final_adder.U$$293/X sky130_fd_sc_hd__a21o_1
XTAP_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$132 U$$678/B1 U$$4/X U$$817/B1 U$$5/X VGND VGND VPWR VPWR U$$133/A sky130_fd_sc_hd__a22o_1
XFILLER_40_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$143 U$$143/A1 U$$165/A2 U$$8/A1 U$$165/B2 VGND VGND VPWR VPWR U$$144/A sky130_fd_sc_hd__a22o_1
XTAP_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$154 U$$154/A U$$176/B VGND VGND VPWR VPWR U$$154/X sky130_fd_sc_hd__xor2_1
XTAP_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_25_1 U$$1121/X U$$1254/X U$$1387/X VGND VGND VPWR VPWR dadda_fa_4_26_0/CIN
+ dadda_fa_4_25_2/A sky130_fd_sc_hd__fa_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$165 U$$28/A1 U$$165/A2 U$$30/A1 U$$165/B2 VGND VGND VPWR VPWR U$$166/A sky130_fd_sc_hd__a22o_1
XTAP_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$176 U$$176/A U$$176/B VGND VGND VPWR VPWR U$$176/X sky130_fd_sc_hd__xor2_1
XFILLER_127_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$187 U$$48/B1 U$$217/A2 U$$598/B1 U$$217/B2 VGND VGND VPWR VPWR U$$188/A sky130_fd_sc_hd__a22o_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$198 U$$198/A U$$218/B VGND VGND VPWR VPWR U$$198/X sky130_fd_sc_hd__xor2_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_18_0 U$$43/X U$$176/X U$$309/X VGND VGND VPWR VPWR dadda_fa_4_19_1/A dadda_fa_4_18_2/A
+ sky130_fd_sc_hd__fa_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_397_ _397_/CLK _397_/D VGND VGND VPWR VPWR _397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1010 U$$2202/B1 VGND VGND VPWR VPWR U$$2065/B1 sky130_fd_sc_hd__buf_4
Xrepeater1021 input86/X VGND VGND VPWR VPWR U$$4450/A1 sky130_fd_sc_hd__buf_6
Xrepeater1032 input84/X VGND VGND VPWR VPWR U$$3348/B1 sky130_fd_sc_hd__buf_6
XFILLER_127_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1043 U$$882/A1 VGND VGND VPWR VPWR U$$2661/B1 sky130_fd_sc_hd__buf_6
Xrepeater1054 U$$4442/A1 VGND VGND VPWR VPWR U$$3207/B1 sky130_fd_sc_hd__buf_6
XFILLER_175_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1065 U$$52/B1 VGND VGND VPWR VPWR U$$54/A1 sky130_fd_sc_hd__buf_6
XFILLER_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_84_5 dadda_fa_2_84_5/A dadda_fa_2_84_5/B dadda_fa_2_84_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_85_2/A dadda_fa_4_84_0/A sky130_fd_sc_hd__fa_2
Xrepeater1076 U$$3612/B1 VGND VGND VPWR VPWR U$$463/A1 sky130_fd_sc_hd__buf_6
XFILLER_99_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1087 U$$50/A1 VGND VGND VPWR VPWR U$$3884/B1 sky130_fd_sc_hd__buf_6
Xrepeater1098 U$$969/A1 VGND VGND VPWR VPWR U$$8/B1 sky130_fd_sc_hd__buf_2
XFILLER_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_77_4 dadda_fa_2_77_4/A dadda_fa_2_77_4/B dadda_fa_2_77_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_1/CIN dadda_fa_3_77_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_100_3 U$$3665/X U$$3798/X U$$3931/X VGND VGND VPWR VPWR dadda_fa_3_101_2/B
+ dadda_fa_3_100_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_693 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_114_1 dadda_fa_5_114_1/A dadda_fa_5_114_1/B dadda_fa_5_114_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_115_0/B dadda_fa_7_114_0/A sky130_fd_sc_hd__fa_1
XFILLER_191_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_107_0 dadda_fa_5_107_0/A dadda_fa_5_107_0/B dadda_fa_5_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_108_0/A dadda_fa_6_107_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_72_3 U$$3210/X U$$3343/X U$$3476/X VGND VGND VPWR VPWR dadda_fa_2_73_1/B
+ dadda_fa_2_72_4/B sky130_fd_sc_hd__fa_1
XFILLER_98_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_65_2 U$$3329/X U$$3462/X U$$3595/X VGND VGND VPWR VPWR dadda_fa_2_66_1/A
+ dadda_fa_2_65_4/A sky130_fd_sc_hd__fa_1
XFILLER_63_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_82_0_1853 VGND VGND VPWR VPWR dadda_fa_1_82_0/A dadda_fa_1_82_0_1853/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_86_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_42_1 dadda_fa_4_42_1/A dadda_fa_4_42_1/B dadda_fa_4_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/B dadda_fa_5_42_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_58_1 U$$1985/X U$$2118/X U$$2251/X VGND VGND VPWR VPWR dadda_fa_2_59_0/CIN
+ dadda_fa_2_58_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_35_0 dadda_fa_4_35_0/A dadda_fa_4_35_0/B dadda_fa_4_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/A dadda_fa_5_35_1/A sky130_fd_sc_hd__fa_1
XFILLER_55_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_320_ _329_/CLK _320_/D VGND VGND VPWR VPWR _320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_251_ _384_/CLK _251_/D VGND VGND VPWR VPWR _251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_182_ _337_/CLK _182_/D VGND VGND VPWR VPWR _182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_87_3 dadda_fa_3_87_3/A dadda_fa_3_87_3/B dadda_fa_3_87_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_88_1/B dadda_fa_4_87_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4403 U$$4403/A U$$4403/B VGND VGND VPWR VPWR U$$4403/X sky130_fd_sc_hd__xor2_1
XFILLER_81_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4414 input67/X U$$4388/X input68/X U$$4426/B2 VGND VGND VPWR VPWR U$$4415/A sky130_fd_sc_hd__a22o_1
XFILLER_78_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_60_1 U$$526/X U$$659/X U$$792/X VGND VGND VPWR VPWR dadda_fa_1_61_6/B
+ dadda_fa_1_60_8/A sky130_fd_sc_hd__fa_1
XFILLER_81_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4425 U$$4425/A U$$4425/B VGND VGND VPWR VPWR U$$4425/X sky130_fd_sc_hd__xor2_1
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4436 U$$4436/A1 U$$4388/X U$$4438/A1 U$$4389/X VGND VGND VPWR VPWR U$$4437/A sky130_fd_sc_hd__a22o_1
XU$$4447 U$$4447/A U$$4447/B VGND VGND VPWR VPWR U$$4447/X sky130_fd_sc_hd__xor2_1
XU$$3702 U$$3836/A U$$3702/B VGND VGND VPWR VPWR U$$3702/X sky130_fd_sc_hd__and2_1
XU$$4458 U$$4458/A1 U$$4388/X U$$4460/A1 U$$4476/B2 VGND VGND VPWR VPWR U$$4459/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3713 U$$3713/A1 U$$3753/A2 U$$3852/A1 U$$3753/B2 VGND VGND VPWR VPWR U$$3714/A
+ sky130_fd_sc_hd__a22o_1
XU$$4469 U$$4469/A U$$4469/B VGND VGND VPWR VPWR U$$4469/X sky130_fd_sc_hd__xor2_1
XTAP_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3724 U$$3724/A U$$3740/B VGND VGND VPWR VPWR U$$3724/X sky130_fd_sc_hd__xor2_1
XTAP_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3735 U$$4420/A1 U$$3739/A2 U$$3737/A1 U$$3739/B2 VGND VGND VPWR VPWR U$$3736/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3746 U$$3746/A U$$3754/B VGND VGND VPWR VPWR U$$3746/X sky130_fd_sc_hd__xor2_1
XFILLER_206_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_554 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3757 input82/X U$$3777/A2 input83/X U$$3777/B2 VGND VGND VPWR VPWR U$$3758/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_109_2 dadda_fa_4_109_2/A dadda_fa_4_109_2/B dadda_fa_4_109_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_110_0/CIN dadda_fa_5_109_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3768 U$$3768/A U$$3774/B VGND VGND VPWR VPWR U$$3768/X sky130_fd_sc_hd__xor2_1
XU$$3779 input94/X U$$3833/A2 input95/X U$$3833/B2 VGND VGND VPWR VPWR U$$3780/A sky130_fd_sc_hd__a22o_1
XTAP_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_82_2 dadda_fa_2_82_2/A dadda_fa_2_82_2/B dadda_fa_2_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/A dadda_fa_3_82_3/A sky130_fd_sc_hd__fa_1
XFILLER_88_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1039 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_75_1 dadda_fa_2_75_1/A dadda_fa_2_75_1/B dadda_fa_2_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_0/CIN dadda_fa_3_75_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_52_0 dadda_fa_5_52_0/A dadda_fa_5_52_0/B dadda_fa_5_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_53_0/A dadda_fa_6_52_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_68_0 dadda_fa_2_68_0/A dadda_fa_2_68_0/B dadda_fa_2_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_0/B dadda_fa_3_68_2/B sky130_fd_sc_hd__fa_1
XFILLER_110_551 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1050 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_97_2 dadda_fa_4_97_2/A dadda_fa_4_97_2/B dadda_fa_4_97_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_98_0/CIN dadda_fa_5_97_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_67_0 dadda_fa_7_67_0/A dadda_fa_7_67_0/B dadda_fa_7_67_0/CIN VGND VGND
+ VPWR VPWR _364_/D _235_/D sky130_fd_sc_hd__fa_1
XFILLER_182_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_70_0 U$$2275/X U$$2408/X U$$2541/X VGND VGND VPWR VPWR dadda_fa_2_71_0/B
+ dadda_fa_2_70_3/B sky130_fd_sc_hd__fa_1
XFILLER_87_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3009 U$$3555/B1 U$$3011/A2 U$$3557/B1 U$$3011/B2 VGND VGND VPWR VPWR U$$3010/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2308 U$$936/B1 U$$2308/A2 U$$2445/B1 U$$2308/B2 VGND VGND VPWR VPWR U$$2309/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2319 U$$2319/A U$$2328/A VGND VGND VPWR VPWR U$$2319/X sky130_fd_sc_hd__xor2_1
XFILLER_28_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1607 U$$98/B1 U$$1607/A2 U$$924/A1 U$$1607/B2 VGND VGND VPWR VPWR U$$1608/A sky130_fd_sc_hd__a22o_1
XFILLER_54_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1618 U$$1618/A U$$1628/B VGND VGND VPWR VPWR U$$1618/X sky130_fd_sc_hd__xor2_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1629 U$$1764/B1 U$$1637/A2 U$$2316/A1 U$$1637/B2 VGND VGND VPWR VPWR U$$1630/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_303_ _304_/CLK _303_/D VGND VGND VPWR VPWR _303_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_234_ _363_/CLK _234_/D VGND VGND VPWR VPWR _234_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_92_1 dadda_fa_3_92_1/A dadda_fa_3_92_1/B dadda_fa_3_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_0/CIN dadda_fa_4_92_2/A sky130_fd_sc_hd__fa_1
XFILLER_109_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_85_0 dadda_fa_3_85_0/A dadda_fa_3_85_0/B dadda_fa_3_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_0/B dadda_fa_4_85_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater507 U$$3132/A2 VGND VGND VPWR VPWR U$$3148/A2 sky130_fd_sc_hd__buf_6
XFILLER_172_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater518 U$$2881/X VGND VGND VPWR VPWR U$$2985/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4200 input100/X U$$4210/A2 U$$4476/A1 U$$4210/B2 VGND VGND VPWR VPWR U$$4201/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater529 U$$2844/A2 VGND VGND VPWR VPWR U$$2810/A2 sky130_fd_sc_hd__buf_6
XU$$4211 U$$4211/A U$$4211/B VGND VGND VPWR VPWR U$$4211/X sky130_fd_sc_hd__xor2_1
XFILLER_66_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4222 U$$4496/A1 U$$4226/A2 U$$4498/A1 U$$4226/B2 VGND VGND VPWR VPWR U$$4223/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4233 U$$4233/A U$$4239/B VGND VGND VPWR VPWR U$$4233/X sky130_fd_sc_hd__xor2_1
XFILLER_133_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4244 U$$4516/B1 U$$4114/X U$$4244/B1 U$$4115/X VGND VGND VPWR VPWR U$$4245/A sky130_fd_sc_hd__a22o_1
XU$$3510 U$$3510/A U$$3510/B VGND VGND VPWR VPWR U$$3510/X sky130_fd_sc_hd__xor2_1
XFILLER_77_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_114_0 U$$4092/X U$$4225/X U$$4358/X VGND VGND VPWR VPWR dadda_fa_5_115_0/A
+ dadda_fa_5_114_1/A sky130_fd_sc_hd__fa_1
XFILLER_19_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4255 U$$4392/A1 U$$4275/A2 U$$4394/A1 U$$4275/B2 VGND VGND VPWR VPWR U$$4256/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_47_5 dadda_fa_2_47_5/A dadda_fa_2_47_5/B dadda_fa_2_47_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_48_2/A dadda_fa_4_47_0/A sky130_fd_sc_hd__fa_1
XFILLER_207_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3521 U$$918/A1 U$$3527/A2 U$$783/A1 U$$3527/B2 VGND VGND VPWR VPWR U$$3522/A sky130_fd_sc_hd__a22o_1
XU$$4266 U$$4266/A U$$4310/B VGND VGND VPWR VPWR U$$4266/X sky130_fd_sc_hd__xor2_1
XFILLER_65_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3532 U$$3532/A U$$3550/B VGND VGND VPWR VPWR U$$3532/X sky130_fd_sc_hd__xor2_1
XFILLER_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4277 input67/X U$$4297/A2 U$$4277/B1 U$$4297/B2 VGND VGND VPWR VPWR U$$4278/A
+ sky130_fd_sc_hd__a22o_1
XU$$3543 U$$3817/A1 U$$3549/A2 U$$3545/A1 U$$3549/B2 VGND VGND VPWR VPWR U$$3544/A
+ sky130_fd_sc_hd__a22o_1
XU$$4288 U$$4288/A U$$4294/B VGND VGND VPWR VPWR U$$4288/X sky130_fd_sc_hd__xor2_1
XFILLER_207_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3554 U$$3554/A U$$3561/A VGND VGND VPWR VPWR U$$3554/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2820 U$$4188/B1 U$$2858/A2 input95/X U$$2858/B2 VGND VGND VPWR VPWR U$$2821/A
+ sky130_fd_sc_hd__a22o_1
XU$$4299 U$$4436/A1 U$$4381/A2 U$$4438/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4300/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3565 U$$3643/B U$$3565/B VGND VGND VPWR VPWR U$$3565/X sky130_fd_sc_hd__and2_1
XU$$3576 U$$3713/A1 U$$3660/A2 U$$3578/A1 U$$3660/B2 VGND VGND VPWR VPWR U$$3577/A
+ sky130_fd_sc_hd__a22o_1
XU$$2831 U$$2831/A U$$2845/B VGND VGND VPWR VPWR U$$2831/X sky130_fd_sc_hd__xor2_1
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2842 U$$2842/A1 U$$2744/X U$$2842/B1 U$$2745/X VGND VGND VPWR VPWR U$$2843/A sky130_fd_sc_hd__a22o_1
XFILLER_34_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3587 U$$3587/A U$$3613/B VGND VGND VPWR VPWR U$$3587/X sky130_fd_sc_hd__xor2_1
XU$$2853 U$$2853/A U$$2876/A VGND VGND VPWR VPWR U$$2853/X sky130_fd_sc_hd__xor2_1
XU$$3598 U$$4420/A1 U$$3636/A2 U$$3737/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3599/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2864 U$$3547/B1 U$$2868/A2 U$$3414/A1 U$$2868/B2 VGND VGND VPWR VPWR U$$2865/A
+ sky130_fd_sc_hd__a22o_1
XU$$2875 U$$2875/A U$$2876/A VGND VGND VPWR VPWR U$$2875/X sky130_fd_sc_hd__xor2_1
XFILLER_179_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2886 U$$2886/A U$$2922/B VGND VGND VPWR VPWR U$$2886/X sky130_fd_sc_hd__xor2_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2897 U$$4404/A1 U$$2919/A2 U$$3447/A1 U$$2919/B2 VGND VGND VPWR VPWR U$$2898/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_191 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$815 final_adder.U$$782/A final_adder.U$$735/X final_adder.U$$703/X
+ VGND VGND VPWR VPWR final_adder.U$$815/X sky130_fd_sc_hd__a21o_2
XFILLER_69_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$837 final_adder.U$$740/X final_adder.U$$805/X final_adder.U$$741/X
+ VGND VGND VPWR VPWR final_adder.U$$837/X sky130_fd_sc_hd__a21o_4
XFILLER_151_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$859 final_adder.U$$762/X final_adder.U$$827/X final_adder.U$$763/X
+ VGND VGND VPWR VPWR final_adder.U$$859/X sky130_fd_sc_hd__a21o_2
XU$$709 U$$709/A1 U$$711/A2 U$$846/B1 U$$711/B2 VGND VGND VPWR VPWR U$$710/A sky130_fd_sc_hd__a22o_1
XFILLER_72_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1609 U$$4494/A1 VGND VGND VPWR VPWR U$$384/A1 sky130_fd_sc_hd__buf_8
XFILLER_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_109_1 U$$3550/X U$$3683/X U$$3816/X VGND VGND VPWR VPWR dadda_fa_4_110_0/CIN
+ dadda_fa_4_109_2/A sky130_fd_sc_hd__fa_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1091 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2105 U$$3749/A1 U$$2113/A2 U$$3749/B1 U$$2113/B2 VGND VGND VPWR VPWR U$$2106/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2116 U$$2116/A U$$2191/A VGND VGND VPWR VPWR U$$2116/X sky130_fd_sc_hd__xor2_1
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2127 U$$894/A1 U$$2169/A2 U$$3499/A1 U$$2169/B2 VGND VGND VPWR VPWR U$$2128/A
+ sky130_fd_sc_hd__a22o_1
XU$$2138 U$$2138/A U$$2170/B VGND VGND VPWR VPWR U$$2138/X sky130_fd_sc_hd__xor2_1
XU$$2149 U$$2834/A1 U$$2149/A2 U$$2425/A1 U$$2149/B2 VGND VGND VPWR VPWR U$$2150/A
+ sky130_fd_sc_hd__a22o_1
XU$$1404 U$$854/B1 U$$1404/A2 U$$719/B1 U$$1404/B2 VGND VGND VPWR VPWR U$$1405/A sky130_fd_sc_hd__a22o_1
XFILLER_27_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1415 U$$1415/A U$$1423/B VGND VGND VPWR VPWR U$$1415/X sky130_fd_sc_hd__xor2_1
XFILLER_188_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1426 U$$328/B1 U$$1462/A2 U$$56/B1 U$$1462/B2 VGND VGND VPWR VPWR U$$1427/A sky130_fd_sc_hd__a22o_1
XFILLER_188_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1437 U$$1437/A U$$1449/B VGND VGND VPWR VPWR U$$1437/X sky130_fd_sc_hd__xor2_1
XFILLER_204_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1448 U$$1448/A1 U$$1448/A2 U$$902/A1 U$$1448/B2 VGND VGND VPWR VPWR U$$1449/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1459 U$$1459/A U$$1459/B VGND VGND VPWR VPWR U$$1459/X sky130_fd_sc_hd__xor2_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_217_ _219_/CLK _217_/D VGND VGND VPWR VPWR _217_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_129_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_974 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_52_3 dadda_fa_2_52_3/A dadda_fa_2_52_3/B dadda_fa_2_52_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/B dadda_fa_3_52_3/B sky130_fd_sc_hd__fa_1
XFILLER_39_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4030 U$$4030/A U$$4036/B VGND VGND VPWR VPWR U$$4030/X sky130_fd_sc_hd__xor2_1
XU$$4041 U$$4176/B1 U$$3977/X U$$4043/A1 U$$3978/X VGND VGND VPWR VPWR U$$4042/A sky130_fd_sc_hd__a22o_1
XU$$4052 U$$4052/A U$$4080/B VGND VGND VPWR VPWR U$$4052/X sky130_fd_sc_hd__xor2_1
XFILLER_211_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4063 input100/X U$$4077/A2 U$$4476/A1 U$$4077/B2 VGND VGND VPWR VPWR U$$4064/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_45_2 input196/X dadda_fa_2_45_2/B dadda_fa_2_45_2/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_46_1/A dadda_fa_3_45_3/A sky130_fd_sc_hd__fa_1
XFILLER_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4074 U$$4074/A U$$4078/B VGND VGND VPWR VPWR U$$4074/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4085 U$$4496/A1 U$$4101/A2 input113/X U$$4101/B2 VGND VGND VPWR VPWR U$$4086/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_22_1 dadda_fa_5_22_1/A dadda_fa_5_22_1/B dadda_fa_5_22_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_23_0/B dadda_fa_7_22_0/A sky130_fd_sc_hd__fa_1
XFILLER_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3340 U$$3612/B1 U$$3348/A2 U$$4027/A1 U$$3346/B2 VGND VGND VPWR VPWR U$$3341/A
+ sky130_fd_sc_hd__a22o_1
XU$$4096 U$$4096/A U$$4100/B VGND VGND VPWR VPWR U$$4096/X sky130_fd_sc_hd__xor2_1
XU$$3351 U$$3351/A U$$3395/B VGND VGND VPWR VPWR U$$3351/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_38_1 U$$1546/X U$$1679/X U$$1812/X VGND VGND VPWR VPWR dadda_fa_3_39_0/CIN
+ dadda_fa_3_38_2/CIN sky130_fd_sc_hd__fa_1
XU$$3362 U$$3908/B1 U$$3378/A2 U$$3775/A1 U$$3378/B2 VGND VGND VPWR VPWR U$$3363/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3373 U$$3373/A U$$3375/B VGND VGND VPWR VPWR U$$3373/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3384 U$$4478/B1 U$$3388/A2 U$$783/A1 U$$3390/B2 VGND VGND VPWR VPWR U$$3385/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_15_0 dadda_fa_5_15_0/A dadda_fa_5_15_0/B dadda_fa_5_15_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_16_0/A dadda_fa_6_15_0/CIN sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_45_clk _385_/CLK VGND VGND VPWR VPWR _387_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_185_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3395 U$$3395/A U$$3395/B VGND VGND VPWR VPWR U$$3395/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2650 U$$2650/A U$$2650/B VGND VGND VPWR VPWR U$$2650/X sky130_fd_sc_hd__xor2_1
XU$$2661 U$$3207/B1 U$$2691/A2 U$$2661/B1 U$$2691/B2 VGND VGND VPWR VPWR U$$2662/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2672 U$$2672/A U$$2680/B VGND VGND VPWR VPWR U$$2672/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2683 U$$4188/B1 U$$2683/A2 U$$2683/B1 U$$2683/B2 VGND VGND VPWR VPWR U$$2684/A
+ sky130_fd_sc_hd__a22o_1
XU$$2694 U$$2694/A U$$2716/B VGND VGND VPWR VPWR U$$2694/X sky130_fd_sc_hd__xor2_1
XFILLER_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1960 U$$3876/B1 U$$1960/A2 U$$864/B1 U$$1960/B2 VGND VGND VPWR VPWR U$$1961/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1971 U$$1971/A U$$1971/B VGND VGND VPWR VPWR U$$1971/X sky130_fd_sc_hd__xor2_1
XU$$1982 input85/X U$$2052/A2 U$$4450/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$1983/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1993 U$$1993/A U$$1993/B VGND VGND VPWR VPWR U$$1993/X sky130_fd_sc_hd__xor2_1
XU$$4405_1779 VGND VGND VPWR VPWR U$$4405_1779/HI U$$4405/B sky130_fd_sc_hd__conb_1
XFILLER_194_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_833 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_941 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_899 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput107 b[48] VGND VGND VPWR VPWR input107/X sky130_fd_sc_hd__buf_6
Xdadda_ha_1_41_3 U$$1286/X U$$1419/X VGND VGND VPWR VPWR dadda_fa_2_42_4/B dadda_fa_3_41_0/A
+ sky130_fd_sc_hd__ha_1
Xinput118 b[58] VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__buf_6
XFILLER_131_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput129 c[0] VGND VGND VPWR VPWR _296_/D sky130_fd_sc_hd__buf_4
XTAP_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$601 final_adder.U$$600/B final_adder.U$$485/X final_adder.U$$477/X
+ VGND VGND VPWR VPWR final_adder.U$$601/X sky130_fd_sc_hd__a21o_1
XTAP_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$612 final_adder.U$$612/A final_adder.U$$612/B VGND VGND VPWR VPWR
+ final_adder.U$$716/A sky130_fd_sc_hd__and2_1
XTAP_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$623 final_adder.U$$614/A final_adder.U$$381/X final_adder.U$$499/X
+ VGND VGND VPWR VPWR final_adder.U$$623/X sky130_fd_sc_hd__a21o_2
XTAP_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$634 final_adder.U$$650/B final_adder.U$$634/B VGND VGND VPWR VPWR
+ final_adder.U$$746/B sky130_fd_sc_hd__and2_1
Xdadda_ha_4_11_1 U$$428/X U$$561/X VGND VGND VPWR VPWR dadda_fa_5_12_0/CIN dadda_ha_4_11_1/SUM
+ sky130_fd_sc_hd__ha_1
XTAP_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$645 final_adder.U$$644/B final_adder.U$$541/X final_adder.U$$525/X
+ VGND VGND VPWR VPWR final_adder.U$$645/X sky130_fd_sc_hd__a21o_1
XFILLER_186_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$656 final_adder.U$$672/B final_adder.U$$656/B VGND VGND VPWR VPWR
+ final_adder.U$$768/B sky130_fd_sc_hd__and2_1
XTAP_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater860 U$$259/B2 VGND VGND VPWR VPWR U$$257/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$667 final_adder.U$$666/B final_adder.U$$563/X final_adder.U$$547/X
+ VGND VGND VPWR VPWR final_adder.U$$667/X sky130_fd_sc_hd__a21o_1
XTAP_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater871 U$$1349/B2 VGND VGND VPWR VPWR U$$1307/B2 sky130_fd_sc_hd__clkbuf_8
XU$$506 U$$506/A U$$528/B VGND VGND VPWR VPWR U$$506/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$678 final_adder.U$$694/B final_adder.U$$678/B VGND VGND VPWR VPWR
+ final_adder.U$$790/B sky130_fd_sc_hd__and2_1
XTAP_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$517 U$$517/A1 U$$521/A2 U$$517/B1 U$$521/B2 VGND VGND VPWR VPWR U$$518/A sky130_fd_sc_hd__a22o_1
XFILLER_29_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater882 U$$1222/B2 VGND VGND VPWR VPWR U$$1190/B2 sky130_fd_sc_hd__buf_8
Xfinal_adder.U$$689 final_adder.U$$688/B final_adder.U$$585/X final_adder.U$$569/X
+ VGND VGND VPWR VPWR final_adder.U$$689/X sky130_fd_sc_hd__a21o_1
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater893 U$$94/B2 VGND VGND VPWR VPWR U$$134/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_40_1 U$$486/X U$$619/X U$$752/X VGND VGND VPWR VPWR dadda_fa_2_41_4/A
+ dadda_fa_2_40_5/B sky130_fd_sc_hd__fa_1
XU$$528 U$$528/A U$$528/B VGND VGND VPWR VPWR U$$528/X sky130_fd_sc_hd__xor2_1
XU$$539 U$$676/A1 U$$415/X U$$676/B1 U$$416/X VGND VGND VPWR VPWR U$$540/A sky130_fd_sc_hd__a22o_1
XFILLER_71_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_983 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_80 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1406 U$$2100/B VGND VGND VPWR VPWR U$$2114/B sky130_fd_sc_hd__buf_6
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1417 U$$2047/B VGND VGND VPWR VPWR U$$2054/A sky130_fd_sc_hd__buf_8
Xrepeater1428 input20/X VGND VGND VPWR VPWR U$$1912/B sky130_fd_sc_hd__buf_4
XFILLER_67_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1439 U$$1628/B VGND VGND VPWR VPWR U$$1620/B sky130_fd_sc_hd__buf_6
XFILLER_125_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_62_2 dadda_fa_3_62_2/A dadda_fa_3_62_2/B dadda_fa_3_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_1/A dadda_fa_4_62_2/B sky130_fd_sc_hd__fa_1
XFILLER_122_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_55_1 dadda_fa_3_55_1/A dadda_fa_3_55_1/B dadda_fa_3_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_0/CIN dadda_fa_4_55_2/A sky130_fd_sc_hd__fa_1
XFILLER_94_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_32_0 dadda_fa_6_32_0/A dadda_fa_6_32_0/B dadda_fa_6_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_33_0/B dadda_fa_7_32_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_208_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_48_0 dadda_fa_3_48_0/A dadda_fa_3_48_0/B dadda_fa_3_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_0/B dadda_fa_4_48_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk _255_/CLK VGND VGND VPWR VPWR _408_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1201 U$$1201/A U$$1205/B VGND VGND VPWR VPWR U$$1201/X sky130_fd_sc_hd__xor2_1
XU$$1212 U$$938/A1 U$$1230/A2 U$$527/B1 U$$1230/B2 VGND VGND VPWR VPWR U$$1213/A sky130_fd_sc_hd__a22o_1
XU$$1223 U$$1223/A U$$1223/B VGND VGND VPWR VPWR U$$1223/X sky130_fd_sc_hd__xor2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1234 input10/X VGND VGND VPWR VPWR U$$1236/B sky130_fd_sc_hd__inv_1
XFILLER_15_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1245 U$$2202/B1 U$$1311/A2 U$$14/A1 U$$1271/B2 VGND VGND VPWR VPWR U$$1246/A sky130_fd_sc_hd__a22o_1
XFILLER_71_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1256 U$$1256/A U$$1270/B VGND VGND VPWR VPWR U$$1256/X sky130_fd_sc_hd__xor2_1
XFILLER_204_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1267 U$$854/B1 U$$1271/A2 U$$719/B1 U$$1271/B2 VGND VGND VPWR VPWR U$$1268/A sky130_fd_sc_hd__a22o_1
XU$$1278 U$$1278/A U$$1286/B VGND VGND VPWR VPWR U$$1278/X sky130_fd_sc_hd__xor2_1
XFILLER_188_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1289 U$$328/B1 U$$1289/A2 U$$58/A1 U$$1291/B2 VGND VGND VPWR VPWR U$$1290/A sky130_fd_sc_hd__a22o_1
XFILLER_206_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_105_0 dadda_fa_7_105_0/A dadda_fa_7_105_0/B dadda_fa_7_105_0/CIN VGND
+ VGND VPWR VPWR _402_/D _273_/D sky130_fd_sc_hd__fa_1
XFILLER_15_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1050 final_adder.U$$228/A final_adder.U$$729/X VGND VGND VPWR VPWR
+ output303/A sky130_fd_sc_hd__xor2_1
XFILLER_8_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1061 final_adder.U$$218/B final_adder.U$$989/X VGND VGND VPWR VPWR
+ output315/A sky130_fd_sc_hd__xor2_1
XFILLER_183_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1072 final_adder.U$$206/A final_adder.U$$819/X VGND VGND VPWR VPWR
+ output327/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1083 final_adder.U$$196/B final_adder.U$$967/X VGND VGND VPWR VPWR
+ output339/A sky130_fd_sc_hd__xor2_1
XFILLER_132_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1094 final_adder.U$$184/A final_adder.U$$893/X VGND VGND VPWR VPWR
+ output352/A sky130_fd_sc_hd__xor2_1
XFILLER_176_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_50_0 U$$3454/B input202/X dadda_fa_2_50_0/CIN VGND VGND VPWR VPWR dadda_fa_3_51_0/B
+ dadda_fa_3_50_2/B sky130_fd_sc_hd__fa_1
XFILLER_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3170 U$$3170/A U$$3264/B VGND VGND VPWR VPWR U$$3170/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_18_clk _380_/CLK VGND VGND VPWR VPWR _246_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3181 input67/X U$$3187/A2 U$$3183/A1 U$$3187/B2 VGND VGND VPWR VPWR U$$3182/A
+ sky130_fd_sc_hd__a22o_1
XU$$3192 U$$3192/A U$$3208/B VGND VGND VPWR VPWR U$$3192/X sky130_fd_sc_hd__xor2_1
XU$$2480 U$$3028/A1 U$$2490/A2 U$$2754/B1 U$$2490/B2 VGND VGND VPWR VPWR U$$2481/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2491 U$$2491/A U$$2491/B VGND VGND VPWR VPWR U$$2491/X sky130_fd_sc_hd__xor2_1
XFILLER_50_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1790 U$$1790/A U$$1820/B VGND VGND VPWR VPWR U$$1790/X sky130_fd_sc_hd__xor2_1
XFILLER_107_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_72_1 dadda_fa_4_72_1/A dadda_fa_4_72_1/B dadda_fa_4_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/B dadda_fa_5_72_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_88_1 U$$2045/X U$$2178/X U$$2311/X VGND VGND VPWR VPWR dadda_fa_2_89_3/CIN
+ dadda_fa_2_88_5/A sky130_fd_sc_hd__fa_1
XFILLER_27_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1064 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_65_0 dadda_fa_4_65_0/A dadda_fa_4_65_0/B dadda_fa_4_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/A dadda_fa_5_65_1/A sky130_fd_sc_hd__fa_1
XFILLER_115_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$420 final_adder.U$$424/B final_adder.U$$420/B VGND VGND VPWR VPWR
+ final_adder.U$$544/B sky130_fd_sc_hd__and2_1
XTAP_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$431 final_adder.U$$430/B final_adder.U$$309/X final_adder.U$$305/X
+ VGND VGND VPWR VPWR final_adder.U$$431/X sky130_fd_sc_hd__a21o_1
XTAP_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$442 final_adder.U$$446/B final_adder.U$$442/B VGND VGND VPWR VPWR
+ final_adder.U$$566/B sky130_fd_sc_hd__and2_1
XTAP_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$453 final_adder.U$$452/B final_adder.U$$331/X final_adder.U$$327/X
+ VGND VGND VPWR VPWR final_adder.U$$453/X sky130_fd_sc_hd__a21o_1
XTAP_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$464 final_adder.U$$468/B final_adder.U$$464/B VGND VGND VPWR VPWR
+ final_adder.U$$588/B sky130_fd_sc_hd__and2_1
XU$$303 U$$303/A U$$379/B VGND VGND VPWR VPWR U$$303/X sky130_fd_sc_hd__xor2_1
XTAP_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$475 final_adder.U$$474/B final_adder.U$$353/X final_adder.U$$349/X
+ VGND VGND VPWR VPWR final_adder.U$$475/X sky130_fd_sc_hd__a21o_1
XFILLER_177_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$314 U$$40/A1 U$$340/A2 U$$42/A1 U$$340/B2 VGND VGND VPWR VPWR U$$315/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$486 final_adder.U$$490/B final_adder.U$$486/B VGND VGND VPWR VPWR
+ final_adder.U$$610/B sky130_fd_sc_hd__and2_1
Xrepeater690 U$$4238/B2 VGND VGND VPWR VPWR U$$4226/B2 sky130_fd_sc_hd__clkbuf_4
XTAP_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$325 U$$325/A U$$351/B VGND VGND VPWR VPWR U$$325/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$497 final_adder.U$$496/B final_adder.U$$375/X final_adder.U$$371/X
+ VGND VGND VPWR VPWR final_adder.U$$497/X sky130_fd_sc_hd__a21o_1
XTAP_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$336 U$$882/B1 U$$340/A2 U$$64/A1 U$$340/B2 VGND VGND VPWR VPWR U$$337/A sky130_fd_sc_hd__a22o_1
XTAP_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$347 U$$347/A U$$367/B VGND VGND VPWR VPWR U$$347/X sky130_fd_sc_hd__xor2_1
XFILLER_199_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$358 U$$630/B1 U$$396/A2 U$$86/A1 U$$396/B2 VGND VGND VPWR VPWR U$$359/A sky130_fd_sc_hd__a22o_1
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_79 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$369 U$$369/A U$$377/B VGND VGND VPWR VPWR U$$369/X sky130_fd_sc_hd__xor2_1
XFILLER_199_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4427_1790 VGND VGND VPWR VPWR U$$4427_1790/HI U$$4427/B sky130_fd_sc_hd__conb_1
XFILLER_158_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1203 input65/X VGND VGND VPWR VPWR U$$3979/B1 sky130_fd_sc_hd__buf_6
XFILLER_193_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1214 U$$492/B VGND VGND VPWR VPWR U$$484/B sky130_fd_sc_hd__buf_6
Xrepeater1225 U$$4382/B VGND VGND VPWR VPWR U$$4384/A sky130_fd_sc_hd__buf_4
Xrepeater1236 U$$4239/B VGND VGND VPWR VPWR U$$4227/B sky130_fd_sc_hd__buf_6
XFILLER_154_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1247 U$$395/B VGND VGND VPWR VPWR U$$367/B sky130_fd_sc_hd__buf_8
Xrepeater1258 U$$3947/B VGND VGND VPWR VPWR U$$3927/B sky130_fd_sc_hd__buf_8
XFILLER_5_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1269 U$$3774/B VGND VGND VPWR VPWR U$$3740/B sky130_fd_sc_hd__buf_8
XFILLER_84_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$828_1843 VGND VGND VPWR VPWR U$$828_1843/HI U$$828/A1 sky130_fd_sc_hd__conb_1
XFILLER_208_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$870 U$$48/A1 U$$872/A2 U$$48/B1 U$$872/B2 VGND VGND VPWR VPWR U$$871/A sky130_fd_sc_hd__a22o_1
XU$$1020 U$$1020/A U$$994/B VGND VGND VPWR VPWR U$$1020/X sky130_fd_sc_hd__xor2_1
XU$$881 U$$881/A U$$883/B VGND VGND VPWR VPWR U$$881/X sky130_fd_sc_hd__xor2_1
XFILLER_211_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$892 U$$892/A1 U$$892/A2 U$$894/A1 U$$892/B2 VGND VGND VPWR VPWR U$$893/A sky130_fd_sc_hd__a22o_1
XFILLER_32_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1031 U$$757/A1 U$$1057/A2 U$$483/B1 U$$1057/B2 VGND VGND VPWR VPWR U$$1032/A sky130_fd_sc_hd__a22o_1
XU$$1042 U$$1042/A U$$968/B VGND VGND VPWR VPWR U$$1042/X sky130_fd_sc_hd__xor2_1
XU$$1053 U$$916/A1 U$$965/A2 U$$916/B1 U$$965/B2 VGND VGND VPWR VPWR U$$1054/A sky130_fd_sc_hd__a22o_1
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1064 U$$1064/A U$$1076/B VGND VGND VPWR VPWR U$$1064/X sky130_fd_sc_hd__xor2_1
XFILLER_92_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1075 U$$938/A1 U$$1083/A2 U$$527/B1 U$$1083/B2 VGND VGND VPWR VPWR U$$1076/A sky130_fd_sc_hd__a22o_1
XU$$1086 U$$1086/A U$$1095/A VGND VGND VPWR VPWR U$$1086/X sky130_fd_sc_hd__xor2_1
XU$$1097 input8/X VGND VGND VPWR VPWR U$$1099/B sky130_fd_sc_hd__inv_1
XFILLER_177_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1042 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_82_0 dadda_fa_5_82_0/A dadda_fa_5_82_0/B dadda_fa_5_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_83_0/A dadda_fa_6_82_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_98_0 dadda_fa_2_98_0/A U$$2464/X U$$2597/X VGND VGND VPWR VPWR dadda_fa_3_99_0/CIN
+ dadda_fa_3_98_2/B sky130_fd_sc_hd__fa_1
XFILLER_145_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_7_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _325_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_74_7 input228/X dadda_fa_1_74_7/B dadda_fa_1_74_7/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_75_2/CIN dadda_fa_2_74_5/CIN sky130_fd_sc_hd__fa_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_67_6 dadda_fa_1_67_6/A dadda_fa_1_67_6/B dadda_fa_1_67_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_2/B dadda_fa_2_67_5/B sky130_fd_sc_hd__fa_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_371 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_94_1 U$$2456/X U$$2589/X VGND VGND VPWR VPWR dadda_fa_2_95_5/CIN dadda_fa_3_94_0/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_7_97_0 dadda_fa_7_97_0/A dadda_fa_7_97_0/B dadda_fa_7_97_0/CIN VGND VGND
+ VPWR VPWR _394_/D _265_/D sky130_fd_sc_hd__fa_1
XFILLER_72_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_112_0 dadda_fa_6_112_0/A dadda_fa_6_112_0/B dadda_fa_6_112_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_113_0/B dadda_fa_7_112_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3906 U$$4043/A1 U$$3840/X U$$4043/B1 U$$3841/X VGND VGND VPWR VPWR U$$3907/A sky130_fd_sc_hd__a22o_1
XTAP_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3917 U$$3917/A U$$3947/B VGND VGND VPWR VPWR U$$3917/X sky130_fd_sc_hd__xor2_1
XTAP_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$250 final_adder.U$$4/SUM final_adder.U$$5/SUM VGND VGND VPWR VPWR
+ final_adder.U$$378/B sky130_fd_sc_hd__and2_1
XU$$3928 U$$4476/A1 U$$3946/A2 U$$4476/B1 U$$3946/B2 VGND VGND VPWR VPWR U$$3929/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$261 final_adder.U$$260/B final_adder.U$$135/X final_adder.U$$133/X
+ VGND VGND VPWR VPWR final_adder.U$$261/X sky130_fd_sc_hd__a21o_1
XU$$3939 U$$3939/A U$$3972/A VGND VGND VPWR VPWR U$$3939/X sky130_fd_sc_hd__xor2_1
XTAP_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$100 U$$98/B1 U$$134/A2 U$$787/A1 U$$134/B2 VGND VGND VPWR VPWR U$$101/A sky130_fd_sc_hd__a22o_1
XFILLER_79_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$272 final_adder.U$$274/B final_adder.U$$272/B VGND VGND VPWR VPWR
+ final_adder.U$$398/B sky130_fd_sc_hd__and2_1
XTAP_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$111 U$$111/A U$$111/B VGND VGND VPWR VPWR U$$111/X sky130_fd_sc_hd__xor2_1
XTAP_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$283 final_adder.U$$282/B final_adder.U$$157/X final_adder.U$$155/X
+ VGND VGND VPWR VPWR final_adder.U$$283/X sky130_fd_sc_hd__a21o_1
XTAP_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_32_3 dadda_fa_3_32_3/A dadda_fa_3_32_3/B dadda_fa_3_32_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_33_1/B dadda_fa_4_32_2/CIN sky130_fd_sc_hd__fa_1
XU$$122 U$$122/A1 U$$122/A2 U$$944/B1 U$$122/B2 VGND VGND VPWR VPWR U$$123/A sky130_fd_sc_hd__a22o_1
XTAP_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$294 final_adder.U$$296/B final_adder.U$$294/B VGND VGND VPWR VPWR
+ final_adder.U$$420/B sky130_fd_sc_hd__and2_1
XTAP_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$133 U$$133/A U$$3/A VGND VGND VPWR VPWR U$$133/X sky130_fd_sc_hd__xor2_1
XU$$144 U$$144/A U$$160/B VGND VGND VPWR VPWR U$$144/X sky130_fd_sc_hd__xor2_1
XTAP_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$155 U$$703/A1 U$$165/A2 U$$20/A1 U$$165/B2 VGND VGND VPWR VPWR U$$156/A sky130_fd_sc_hd__a22o_1
XTAP_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$166 U$$166/A U$$184/B VGND VGND VPWR VPWR U$$166/X sky130_fd_sc_hd__xor2_1
XTAP_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_25_2 U$$1520/X U$$1653/X input174/X VGND VGND VPWR VPWR dadda_fa_4_26_1/A
+ dadda_fa_4_25_2/B sky130_fd_sc_hd__fa_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$177 U$$40/A1 U$$209/A2 U$$179/A1 U$$209/B2 VGND VGND VPWR VPWR U$$178/A sky130_fd_sc_hd__a22o_1
XFILLER_73_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$188 U$$188/A U$$218/B VGND VGND VPWR VPWR U$$188/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_18_1 U$$442/X U$$575/X U$$708/X VGND VGND VPWR VPWR dadda_fa_4_19_1/B
+ dadda_fa_4_18_2/B sky130_fd_sc_hd__fa_1
XU$$199 U$$882/B1 U$$217/A2 U$$64/A1 U$$217/B2 VGND VGND VPWR VPWR U$$200/A sky130_fd_sc_hd__a22o_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_942 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_396_ _399_/CLK _396_/D VGND VGND VPWR VPWR _396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1000 U$$342/A1 VGND VGND VPWR VPWR U$$68/A1 sky130_fd_sc_hd__buf_4
XFILLER_182_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1011 U$$3300/A1 VGND VGND VPWR VPWR U$$2202/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_127_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1022 U$$4311/B1 VGND VGND VPWR VPWR U$$4176/A1 sky130_fd_sc_hd__buf_6
Xrepeater1033 U$$610/A1 VGND VGND VPWR VPWR U$$882/B1 sky130_fd_sc_hd__buf_4
Xrepeater1044 U$$3485/A1 VGND VGND VPWR VPWR U$$882/A1 sky130_fd_sc_hd__buf_6
XFILLER_86_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1055 U$$4442/A1 VGND VGND VPWR VPWR U$$4440/B1 sky130_fd_sc_hd__buf_6
Xrepeater1066 U$$3614/B1 VGND VGND VPWR VPWR U$$52/B1 sky130_fd_sc_hd__buf_8
XFILLER_175_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1077 U$$4162/A1 VGND VGND VPWR VPWR U$$3612/B1 sky130_fd_sc_hd__buf_6
XFILLER_142_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1088 input78/X VGND VGND VPWR VPWR U$$4434/A1 sky130_fd_sc_hd__buf_6
XFILLER_141_357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1099 U$$2202/A1 VGND VGND VPWR VPWR U$$969/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_77_5 dadda_fa_2_77_5/A dadda_fa_2_77_5/B dadda_fa_2_77_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_78_2/A dadda_fa_4_77_0/A sky130_fd_sc_hd__fa_2
XFILLER_96_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_934 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_438 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_107_1 dadda_fa_5_107_1/A dadda_fa_5_107_1/B dadda_fa_5_107_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_108_0/B dadda_fa_7_107_0/A sky130_fd_sc_hd__fa_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_72_4 U$$3609/X U$$3742/X U$$3875/X VGND VGND VPWR VPWR dadda_fa_2_73_1/CIN
+ dadda_fa_2_72_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_98_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_65_3 U$$3728/X U$$3861/X U$$3994/X VGND VGND VPWR VPWR dadda_fa_2_66_1/B
+ dadda_fa_2_65_4/B sky130_fd_sc_hd__fa_1
XFILLER_63_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_42_2 dadda_fa_4_42_2/A dadda_fa_4_42_2/B dadda_fa_4_42_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_43_0/CIN dadda_fa_5_42_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_2 U$$2384/X U$$2517/X U$$2650/X VGND VGND VPWR VPWR dadda_fa_2_59_1/A
+ dadda_fa_2_58_4/A sky130_fd_sc_hd__fa_1
XFILLER_27_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_35_1 dadda_fa_4_35_1/A dadda_fa_4_35_1/B dadda_fa_4_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/B dadda_fa_5_35_1/B sky130_fd_sc_hd__fa_1
XFILLER_39_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_12_0 dadda_fa_7_12_0/A dadda_fa_7_12_0/B dadda_fa_7_12_0/CIN VGND VGND
+ VPWR VPWR _309_/D _180_/D sky130_fd_sc_hd__fa_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_28_0 dadda_fa_4_28_0/A dadda_fa_4_28_0/B dadda_fa_4_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/A dadda_fa_5_28_1/A sky130_fd_sc_hd__fa_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_250_ _384_/CLK _250_/D VGND VGND VPWR VPWR _250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_181_ _342_/CLK _181_/D VGND VGND VPWR VPWR _181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_0_61_4 U$$1725/X U$$1858/X VGND VGND VPWR VPWR dadda_fa_1_62_7/A dadda_fa_2_61_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_151_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4404 U$$4404/A1 U$$4388/X U$$4406/A1 U$$4430/B2 VGND VGND VPWR VPWR U$$4405/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4415 U$$4415/A U$$4415/B VGND VGND VPWR VPWR U$$4415/X sky130_fd_sc_hd__xor2_1
XFILLER_65_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_60_2 U$$925/X U$$1058/X U$$1191/X VGND VGND VPWR VPWR dadda_fa_1_61_6/CIN
+ dadda_fa_1_60_8/B sky130_fd_sc_hd__fa_1
XU$$4426 U$$4426/A1 U$$4388/X U$$4428/A1 U$$4426/B2 VGND VGND VPWR VPWR U$$4427/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4437 U$$4437/A U$$4437/B VGND VGND VPWR VPWR U$$4437/X sky130_fd_sc_hd__xor2_1
XTAP_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3703 U$$3701/Y input50/X input49/X U$$3702/X U$$3699/Y VGND VGND VPWR VPWR U$$3703/X
+ sky130_fd_sc_hd__a32o_4
XTAP_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4448 input85/X U$$4388/X input86/X U$$4498/B2 VGND VGND VPWR VPWR U$$4449/A sky130_fd_sc_hd__a22o_1
XU$$4459 U$$4459/A U$$4459/B VGND VGND VPWR VPWR U$$4459/X sky130_fd_sc_hd__xor2_1
XTAP_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3714 U$$3714/A U$$3754/B VGND VGND VPWR VPWR U$$3714/X sky130_fd_sc_hd__xor2_1
XU$$3725 U$$4408/B1 U$$3739/A2 U$$4275/A1 U$$3739/B2 VGND VGND VPWR VPWR U$$3726/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3736 U$$3736/A U$$3740/B VGND VGND VPWR VPWR U$$3736/X sky130_fd_sc_hd__xor2_1
XTAP_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3747 U$$3747/A1 U$$3753/A2 U$$50/A1 U$$3753/B2 VGND VGND VPWR VPWR U$$3748/A sky130_fd_sc_hd__a22o_1
XTAP_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_0 U$$1929/X U$$2062/X U$$2094/B VGND VGND VPWR VPWR dadda_fa_4_31_0/B
+ dadda_fa_4_30_1/CIN sky130_fd_sc_hd__fa_1
XU$$3758 U$$3758/A U$$3778/B VGND VGND VPWR VPWR U$$3758/X sky130_fd_sc_hd__xor2_1
XFILLER_205_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3769 U$$4043/A1 U$$3773/A2 U$$4043/B1 U$$3773/B2 VGND VGND VPWR VPWR U$$3770/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_379_ _379_/CLK _379_/D VGND VGND VPWR VPWR _379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_82_3 dadda_fa_2_82_3/A dadda_fa_2_82_3/B dadda_fa_2_82_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/B dadda_fa_3_82_3/B sky130_fd_sc_hd__fa_1
XFILLER_115_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_75_2 dadda_fa_2_75_2/A dadda_fa_2_75_2/B dadda_fa_2_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/A dadda_fa_3_75_3/A sky130_fd_sc_hd__fa_1
XFILLER_141_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_52_1 dadda_fa_5_52_1/A dadda_fa_5_52_1/B dadda_fa_5_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_53_0/B dadda_fa_7_52_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_68_1 dadda_fa_2_68_1/A dadda_fa_2_68_1/B dadda_fa_2_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_0/CIN dadda_fa_3_68_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_45_0 dadda_fa_5_45_0/A dadda_fa_5_45_0/B dadda_fa_5_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_46_0/A dadda_fa_6_45_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_70_1 U$$2674/X U$$2807/X U$$2940/X VGND VGND VPWR VPWR dadda_fa_2_71_0/CIN
+ dadda_fa_2_70_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_0 U$$2394/X U$$2527/X U$$2660/X VGND VGND VPWR VPWR dadda_fa_2_64_0/B
+ dadda_fa_2_63_3/B sky130_fd_sc_hd__fa_1
XFILLER_75_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2309 U$$2309/A U$$2309/B VGND VGND VPWR VPWR U$$2309/X sky130_fd_sc_hd__xor2_1
XFILLER_76_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1608 U$$1608/A U$$1608/B VGND VGND VPWR VPWR U$$1608/X sky130_fd_sc_hd__xor2_1
XU$$1619 U$$521/B1 U$$1621/A2 U$$660/B1 U$$1621/B2 VGND VGND VPWR VPWR U$$1620/A sky130_fd_sc_hd__a22o_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ _304_/CLK _302_/D VGND VGND VPWR VPWR _302_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_233_ _363_/CLK _233_/D VGND VGND VPWR VPWR _233_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_204_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_92_2 dadda_fa_3_92_2/A dadda_fa_3_92_2/B dadda_fa_3_92_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_1/A dadda_fa_4_92_2/B sky130_fd_sc_hd__fa_1
XFILLER_7_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_85_1 dadda_fa_3_85_1/A dadda_fa_3_85_1/B dadda_fa_3_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_0/CIN dadda_fa_4_85_2/A sky130_fd_sc_hd__fa_1
XFILLER_83_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_62_0 dadda_fa_6_62_0/A dadda_fa_6_62_0/B dadda_fa_6_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_63_0/B dadda_fa_7_62_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_78_0 dadda_fa_3_78_0/A dadda_fa_3_78_0/B dadda_fa_3_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_0/B dadda_fa_4_78_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_52_0 U$$111/X U$$244/X VGND VGND VPWR VPWR dadda_fa_1_53_8/CIN dadda_fa_2_52_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_112_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater508 U$$3118/A2 VGND VGND VPWR VPWR U$$3132/A2 sky130_fd_sc_hd__buf_4
XU$$4201 U$$4201/A U$$4211/B VGND VGND VPWR VPWR U$$4201/X sky130_fd_sc_hd__xor2_1
Xrepeater519 U$$396/A2 VGND VGND VPWR VPWR U$$350/A2 sky130_fd_sc_hd__buf_6
XU$$4212 U$$4484/B1 U$$4226/A2 U$$789/A1 U$$4226/B2 VGND VGND VPWR VPWR U$$4213/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4223 U$$4223/A U$$4227/B VGND VGND VPWR VPWR U$$4223/X sky130_fd_sc_hd__xor2_1
XFILLER_77_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4234 U$$4369/B1 U$$4238/A2 U$$4236/A1 U$$4238/B2 VGND VGND VPWR VPWR U$$4235/A
+ sky130_fd_sc_hd__a22o_1
XU$$3500 U$$3500/A U$$3504/B VGND VGND VPWR VPWR U$$3500/X sky130_fd_sc_hd__xor2_1
XU$$4245 U$$4245/A U$$4246/A VGND VGND VPWR VPWR U$$4245/X sky130_fd_sc_hd__xor2_1
XFILLER_19_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4256 U$$4256/A U$$4278/B VGND VGND VPWR VPWR U$$4256/X sky130_fd_sc_hd__xor2_1
XU$$3511 U$$3511/A1 U$$3517/A2 U$$3648/B1 U$$3517/B2 VGND VGND VPWR VPWR U$$3512/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_114_1 U$$4491/X input145/X dadda_fa_4_114_1/CIN VGND VGND VPWR VPWR dadda_fa_5_115_0/B
+ dadda_fa_5_114_1/B sky130_fd_sc_hd__fa_1
XU$$3522 U$$3522/A U$$3528/B VGND VGND VPWR VPWR U$$3522/X sky130_fd_sc_hd__xor2_1
XU$$4267 U$$4402/B1 U$$4297/A2 U$$4406/A1 U$$4297/B2 VGND VGND VPWR VPWR U$$4268/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3533 U$$3944/A1 U$$3549/A2 U$$3944/B1 U$$3549/B2 VGND VGND VPWR VPWR U$$3534/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4278 U$$4278/A U$$4278/B VGND VGND VPWR VPWR U$$4278/X sky130_fd_sc_hd__xor2_1
XU$$3544 U$$3544/A U$$3550/B VGND VGND VPWR VPWR U$$3544/X sky130_fd_sc_hd__xor2_1
XFILLER_81_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4289 U$$4289/A1 U$$4251/X input74/X U$$4252/X VGND VGND VPWR VPWR U$$4290/A sky130_fd_sc_hd__a22o_1
XU$$3555 U$$4240/A1 U$$3559/A2 U$$3555/B1 U$$3559/B2 VGND VGND VPWR VPWR U$$3556/A
+ sky130_fd_sc_hd__a22o_1
XU$$2810 U$$4178/B1 U$$2810/A2 U$$2810/B1 U$$2810/B2 VGND VGND VPWR VPWR U$$2811/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_107_0 dadda_fa_4_107_0/A dadda_fa_4_107_0/B dadda_fa_4_107_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/A dadda_fa_5_107_1/A sky130_fd_sc_hd__fa_1
XU$$2821 U$$2821/A U$$2859/B VGND VGND VPWR VPWR U$$2821/X sky130_fd_sc_hd__xor2_1
XFILLER_65_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3566 U$$3564/Y input48/X input47/X U$$3565/X U$$3562/Y VGND VGND VPWR VPWR U$$3566/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_92_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3577 U$$3577/A U$$3665/B VGND VGND VPWR VPWR U$$3577/X sky130_fd_sc_hd__xor2_1
XU$$2832 U$$3243/A1 U$$2844/A2 U$$3245/A1 U$$2844/B2 VGND VGND VPWR VPWR U$$2833/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2843 U$$2843/A U$$2845/B VGND VGND VPWR VPWR U$$2843/X sky130_fd_sc_hd__xor2_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_806 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3588 U$$4408/B1 U$$3606/A2 U$$4275/A1 U$$3606/B2 VGND VGND VPWR VPWR U$$3589/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2854 U$$660/B1 U$$2858/A2 U$$4361/B1 U$$2858/B2 VGND VGND VPWR VPWR U$$2855/A
+ sky130_fd_sc_hd__a22o_1
XU$$3599 U$$3599/A U$$3637/B VGND VGND VPWR VPWR U$$3599/X sky130_fd_sc_hd__xor2_1
XU$$2865 U$$2865/A U$$2869/B VGND VGND VPWR VPWR U$$2865/X sky130_fd_sc_hd__xor2_1
XU$$2876 U$$2876/A VGND VGND VPWR VPWR U$$2876/Y sky130_fd_sc_hd__inv_1
XFILLER_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2887 U$$3159/B1 U$$2921/A2 U$$3026/A1 U$$2921/B2 VGND VGND VPWR VPWR U$$2888/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_170 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2898 U$$2898/A U$$2920/B VGND VGND VPWR VPWR U$$2898/X sky130_fd_sc_hd__xor2_1
XANTENNA_181 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_80_0 input235/X dadda_fa_2_80_0/B dadda_fa_2_80_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_81_0/B dadda_fa_3_80_2/B sky130_fd_sc_hd__fa_1
XFILLER_143_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_506 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_50_8 U$$3299/X U$$3432/X VGND VGND VPWR VPWR dadda_fa_2_51_3/A dadda_fa_3_50_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_143_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$805 final_adder.U$$772/A final_adder.U$$725/X final_adder.U$$693/X
+ VGND VGND VPWR VPWR final_adder.U$$805/X sky130_fd_sc_hd__a21o_1
XFILLER_5_1218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$827 final_adder.U$$794/A final_adder.U$$503/X final_adder.U$$715/X
+ VGND VGND VPWR VPWR final_adder.U$$827/X sky130_fd_sc_hd__a21o_1
XFILLER_68_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$849 final_adder.U$$752/X final_adder.U$$817/X final_adder.U$$753/X
+ VGND VGND VPWR VPWR final_adder.U$$849/X sky130_fd_sc_hd__a21o_2
XFILLER_57_959 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_812 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_95_0 dadda_fa_4_95_0/A dadda_fa_4_95_0/B dadda_fa_4_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/A dadda_fa_5_95_1/A sky130_fd_sc_hd__fa_1
XFILLER_137_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_109_2 U$$3949/X U$$4082/X U$$4215/X VGND VGND VPWR VPWR dadda_fa_4_110_1/A
+ dadda_fa_4_109_2/B sky130_fd_sc_hd__fa_1
XFILLER_161_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput380 output380/A VGND VGND VPWR VPWR o[96] sky130_fd_sc_hd__buf_2
XFILLER_86_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$965_1845 VGND VGND VPWR VPWR U$$965_1845/HI U$$965/A1 sky130_fd_sc_hd__conb_1
XFILLER_120_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4463_1808 VGND VGND VPWR VPWR U$$4463_1808/HI U$$4463/B sky130_fd_sc_hd__conb_1
XU$$2106 U$$2106/A U$$2114/B VGND VGND VPWR VPWR U$$2106/X sky130_fd_sc_hd__xor2_1
XFILLER_56_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2117 U$$3348/B1 U$$2189/A2 U$$3213/B1 U$$2189/B2 VGND VGND VPWR VPWR U$$2118/A
+ sky130_fd_sc_hd__a22o_1
XU$$2128 U$$2128/A U$$2170/B VGND VGND VPWR VPWR U$$2128/X sky130_fd_sc_hd__xor2_1
XFILLER_76_1011 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2139 U$$3235/A1 U$$2149/A2 U$$2415/A1 U$$2149/B2 VGND VGND VPWR VPWR U$$2140/A
+ sky130_fd_sc_hd__a22o_1
XU$$1405 U$$1405/A U$$1405/B VGND VGND VPWR VPWR U$$1405/X sky130_fd_sc_hd__xor2_1
XFILLER_16_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1416 U$$594/A1 U$$1422/A2 U$$594/B1 U$$1422/B2 VGND VGND VPWR VPWR U$$1417/A sky130_fd_sc_hd__a22o_1
XFILLER_27_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1427 U$$1427/A U$$1459/B VGND VGND VPWR VPWR U$$1427/X sky130_fd_sc_hd__xor2_1
XFILLER_71_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1438 U$$342/A1 U$$1448/A2 U$$1714/A1 U$$1448/B2 VGND VGND VPWR VPWR U$$1439/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1449 U$$1449/A U$$1449/B VGND VGND VPWR VPWR U$$1449/X sky130_fd_sc_hd__xor2_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_216_ _345_/CLK _216_/D VGND VGND VPWR VPWR _216_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_986 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_52_4 dadda_fa_2_52_4/A dadda_fa_2_52_4/B dadda_fa_2_52_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_1/CIN dadda_fa_3_52_3/CIN sky130_fd_sc_hd__fa_1
XU$$4020 U$$4020/A U$$4100/B VGND VGND VPWR VPWR U$$4020/X sky130_fd_sc_hd__xor2_1
XFILLER_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4031 U$$4442/A1 U$$4035/A2 U$$4442/B1 U$$4035/B2 VGND VGND VPWR VPWR U$$4032/A
+ sky130_fd_sc_hd__a22o_1
XU$$4042 U$$4042/A U$$4109/A VGND VGND VPWR VPWR U$$4042/X sky130_fd_sc_hd__xor2_1
XU$$4053 U$$4188/B1 U$$4079/A2 input95/X U$$4079/B2 VGND VGND VPWR VPWR U$$4054/A
+ sky130_fd_sc_hd__a22o_1
XU$$4064 U$$4064/A U$$4078/B VGND VGND VPWR VPWR U$$4064/X sky130_fd_sc_hd__xor2_1
XFILLER_19_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_45_3 dadda_fa_2_45_3/A dadda_fa_2_45_3/B dadda_fa_2_45_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_1/B dadda_fa_3_45_3/B sky130_fd_sc_hd__fa_1
XFILLER_65_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4075 U$$4210/B1 U$$4077/A2 U$$4488/A1 U$$4077/B2 VGND VGND VPWR VPWR U$$4076/A
+ sky130_fd_sc_hd__a22o_1
XU$$3330 U$$4426/A1 U$$3374/A2 U$$4428/A1 U$$3374/B2 VGND VGND VPWR VPWR U$$3331/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4086 U$$4086/A U$$4110/A VGND VGND VPWR VPWR U$$4086/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3341 U$$3341/A U$$3349/B VGND VGND VPWR VPWR U$$3341/X sky130_fd_sc_hd__xor2_1
XU$$3352 U$$3352/A1 U$$3388/A2 input86/X U$$3390/B2 VGND VGND VPWR VPWR U$$3353/A
+ sky130_fd_sc_hd__a22o_1
XU$$4097 U$$4508/A1 U$$4101/A2 U$$4510/A1 U$$4101/B2 VGND VGND VPWR VPWR U$$4098/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_38_2 U$$1945/X U$$2078/X U$$2211/X VGND VGND VPWR VPWR dadda_fa_3_39_1/A
+ dadda_fa_3_38_3/A sky130_fd_sc_hd__fa_1
XU$$3363 U$$3363/A U$$3425/A VGND VGND VPWR VPWR U$$3363/X sky130_fd_sc_hd__xor2_1
XU$$3374 U$$3511/A1 U$$3374/A2 U$$3376/A1 U$$3374/B2 VGND VGND VPWR VPWR U$$3375/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2640 U$$2640/A U$$2650/B VGND VGND VPWR VPWR U$$2640/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_15_1 dadda_fa_5_15_1/A dadda_fa_5_15_1/B dadda_fa_5_15_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_16_0/B dadda_fa_7_15_0/A sky130_fd_sc_hd__fa_1
XU$$3385 U$$3385/A U$$3389/B VGND VGND VPWR VPWR U$$3385/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3396 U$$3944/A1 U$$3416/A2 U$$3944/B1 U$$3416/B2 VGND VGND VPWR VPWR U$$3397/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2651 U$$3747/A1 U$$2653/A2 U$$2925/B1 U$$2653/B2 VGND VGND VPWR VPWR U$$2652/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2662 U$$2662/A U$$2680/B VGND VGND VPWR VPWR U$$2662/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2673 U$$2808/B1 U$$2691/A2 U$$2810/B1 U$$2691/B2 VGND VGND VPWR VPWR U$$2674/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2684 U$$2684/A U$$2736/B VGND VGND VPWR VPWR U$$2684/X sky130_fd_sc_hd__xor2_1
XU$$1950 U$$3594/A1 U$$1960/A2 U$$993/A1 U$$1960/B2 VGND VGND VPWR VPWR U$$1951/A
+ sky130_fd_sc_hd__a22o_1
XU$$2695 U$$3517/A1 U$$2711/A2 U$$3245/A1 U$$2711/B2 VGND VGND VPWR VPWR U$$2696/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1961 U$$1961/A U$$2009/B VGND VGND VPWR VPWR U$$1961/X sky130_fd_sc_hd__xor2_1
XFILLER_167_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1972 U$$3614/B1 U$$2016/A2 U$$3481/A1 U$$2016/B2 VGND VGND VPWR VPWR U$$1973/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1983 U$$1983/A U$$2054/A VGND VGND VPWR VPWR U$$1983/X sky130_fd_sc_hd__xor2_1
XU$$1994 U$$759/B1 U$$2040/A2 U$$763/A1 U$$2040/B2 VGND VGND VPWR VPWR U$$1995/A sky130_fd_sc_hd__a22o_1
XFILLER_31_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput108 b[49] VGND VGND VPWR VPWR input108/X sky130_fd_sc_hd__buf_6
Xinput119 b[59] VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__buf_6
XFILLER_131_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$602 final_adder.U$$610/B final_adder.U$$602/B VGND VGND VPWR VPWR
+ final_adder.U$$706/A sky130_fd_sc_hd__and2_1
XTAP_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$613 final_adder.U$$612/B final_adder.U$$497/X final_adder.U$$489/X
+ VGND VGND VPWR VPWR final_adder.U$$613/X sky130_fd_sc_hd__a21o_1
XFILLER_9_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$635 final_adder.U$$634/B final_adder.U$$531/X final_adder.U$$515/X
+ VGND VGND VPWR VPWR final_adder.U$$635/X sky130_fd_sc_hd__a21o_1
XTAP_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$646 final_adder.U$$662/B final_adder.U$$646/B VGND VGND VPWR VPWR
+ final_adder.U$$758/B sky130_fd_sc_hd__and2_1
XTAP_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater850 U$$1557/B2 VGND VGND VPWR VPWR U$$1545/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$657 final_adder.U$$656/B final_adder.U$$553/X final_adder.U$$537/X
+ VGND VGND VPWR VPWR final_adder.U$$657/X sky130_fd_sc_hd__a21o_1
XTAP_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater861 U$$142/X VGND VGND VPWR VPWR U$$259/B2 sky130_fd_sc_hd__buf_4
XFILLER_110_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$668 final_adder.U$$684/B final_adder.U$$668/B VGND VGND VPWR VPWR
+ final_adder.U$$780/B sky130_fd_sc_hd__and2_1
XTAP_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$507 U$$916/B1 U$$521/A2 U$$920/A1 U$$521/B2 VGND VGND VPWR VPWR U$$508/A sky130_fd_sc_hd__a22o_1
XFILLER_57_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater872 U$$1349/B2 VGND VGND VPWR VPWR U$$1355/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$679 final_adder.U$$678/B final_adder.U$$575/X final_adder.U$$559/X
+ VGND VGND VPWR VPWR final_adder.U$$679/X sky130_fd_sc_hd__a21o_1
XU$$518 U$$518/A U$$528/B VGND VGND VPWR VPWR U$$518/X sky130_fd_sc_hd__xor2_1
XFILLER_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater883 U$$1101/X VGND VGND VPWR VPWR U$$1222/B2 sky130_fd_sc_hd__buf_6
Xrepeater894 U$$5/X VGND VGND VPWR VPWR U$$94/B2 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_1_40_2 U$$885/X U$$1018/X U$$1151/X VGND VGND VPWR VPWR dadda_fa_2_41_4/B
+ dadda_fa_2_40_5/CIN sky130_fd_sc_hd__fa_1
XU$$529 U$$940/A1 U$$537/A2 U$$940/B1 U$$537/B2 VGND VGND VPWR VPWR U$$530/A sky130_fd_sc_hd__a22o_1
XFILLER_38_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_1058 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$90 U$$90/A1 U$$94/A2 U$$92/A1 U$$94/B2 VGND VGND VPWR VPWR U$$91/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_10_0 U$$27/X U$$160/X U$$293/X VGND VGND VPWR VPWR dadda_fa_5_11_0/CIN
+ dadda_fa_5_10_1/B sky130_fd_sc_hd__fa_1
XFILLER_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_70 _342_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_81 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_92 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1407 U$$2150/B VGND VGND VPWR VPWR U$$2100/B sky130_fd_sc_hd__buf_8
XFILLER_125_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_114_0 dadda_fa_3_114_0/A U$$3560/X U$$3693/X VGND VGND VPWR VPWR dadda_fa_4_115_2/A
+ dadda_fa_4_114_2/B sky130_fd_sc_hd__fa_1
Xrepeater1418 U$$2047/B VGND VGND VPWR VPWR U$$2037/B sky130_fd_sc_hd__buf_8
Xrepeater1429 U$$1739/B VGND VGND VPWR VPWR U$$1689/B sky130_fd_sc_hd__buf_6
XFILLER_125_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_62_3 dadda_fa_3_62_3/A dadda_fa_3_62_3/B dadda_fa_3_62_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_63_1/B dadda_fa_4_62_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_121_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_55_2 dadda_fa_3_55_2/A dadda_fa_3_55_2/B dadda_fa_3_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_1/A dadda_fa_4_55_2/B sky130_fd_sc_hd__fa_1
XFILLER_47_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_48_1 dadda_fa_3_48_1/A dadda_fa_3_48_1/B dadda_fa_3_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_0/CIN dadda_fa_4_48_2/A sky130_fd_sc_hd__fa_1
XFILLER_47_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_25_0 dadda_fa_6_25_0/A dadda_fa_6_25_0/B dadda_fa_6_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_26_0/B dadda_fa_7_25_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_169_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1202 U$$2709/A1 U$$1204/A2 U$$2709/B1 U$$1204/B2 VGND VGND VPWR VPWR U$$1203/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1213 U$$1213/A U$$1232/A VGND VGND VPWR VPWR U$$1213/X sky130_fd_sc_hd__xor2_1
XFILLER_16_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1224 U$$2318/B1 U$$1230/A2 U$$952/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1225/A
+ sky130_fd_sc_hd__a22o_1
XU$$1235 U$$1338/B VGND VGND VPWR VPWR U$$1235/Y sky130_fd_sc_hd__inv_1
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1246 U$$1246/A U$$1272/B VGND VGND VPWR VPWR U$$1246/X sky130_fd_sc_hd__xor2_1
XFILLER_15_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1257 U$$1666/B1 U$$1289/A2 U$$985/A1 U$$1281/B2 VGND VGND VPWR VPWR U$$1258/A
+ sky130_fd_sc_hd__a22o_1
XU$$1268 U$$1268/A U$$1270/B VGND VGND VPWR VPWR U$$1268/X sky130_fd_sc_hd__xor2_1
XU$$1279 U$$731/A1 U$$1323/A2 U$$733/A1 U$$1307/B2 VGND VGND VPWR VPWR U$$1280/A sky130_fd_sc_hd__a22o_1
XFILLER_203_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1040 final_adder.U$$238/A final_adder.U$$619/X VGND VGND VPWR VPWR
+ output292/A sky130_fd_sc_hd__xor2_1
XFILLER_172_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1051 final_adder.U$$228/B final_adder.U$$999/X VGND VGND VPWR VPWR
+ output304/A sky130_fd_sc_hd__xor2_1
XFILLER_176_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1062 final_adder.U$$216/A final_adder.U$$829/X VGND VGND VPWR VPWR
+ output316/A sky130_fd_sc_hd__xor2_1
XFILLER_176_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1073 final_adder.U$$206/B final_adder.U$$977/X VGND VGND VPWR VPWR
+ output328/A sky130_fd_sc_hd__xor2_1
XFILLER_183_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1084 final_adder.U$$194/A final_adder.U$$807/X VGND VGND VPWR VPWR
+ output341/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1095 final_adder.U$$184/B final_adder.U$$955/X VGND VGND VPWR VPWR
+ output353/A sky130_fd_sc_hd__xor2_1
XFILLER_171_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_731 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_50_1 dadda_fa_2_50_1/A dadda_fa_2_50_1/B dadda_fa_2_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_0/CIN dadda_fa_3_50_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_43_0 U$$1955/X U$$2088/X U$$2221/X VGND VGND VPWR VPWR dadda_fa_3_44_0/B
+ dadda_fa_3_43_2/B sky130_fd_sc_hd__fa_1
XFILLER_54_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3160 U$$3160/A U$$3208/B VGND VGND VPWR VPWR U$$3160/X sky130_fd_sc_hd__xor2_1
XU$$3171 U$$431/A1 U$$3263/A2 U$$842/B1 U$$3263/B2 VGND VGND VPWR VPWR U$$3172/A sky130_fd_sc_hd__a22o_1
XFILLER_53_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3182 U$$3182/A U$$3188/B VGND VGND VPWR VPWR U$$3182/X sky130_fd_sc_hd__xor2_1
XU$$3193 U$$727/A1 U$$3207/A2 U$$727/B1 U$$3207/B2 VGND VGND VPWR VPWR U$$3194/A sky130_fd_sc_hd__a22o_1
XFILLER_59_1072 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2470 U$$2468/Y input30/X U$$2466/A U$$2469/X U$$2466/Y VGND VGND VPWR VPWR U$$2470/X
+ sky130_fd_sc_hd__a32o_4
XU$$2481 U$$2481/A U$$2491/B VGND VGND VPWR VPWR U$$2481/X sky130_fd_sc_hd__xor2_1
XFILLER_21_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2492 U$$2492/A1 U$$2524/A2 U$$3453/A1 U$$2524/B2 VGND VGND VPWR VPWR U$$2493/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1780 U$$1780/A VGND VGND VPWR VPWR U$$1780/Y sky130_fd_sc_hd__inv_1
XU$$1791 U$$2063/B1 U$$1819/A2 U$$2065/B1 U$$1819/B2 VGND VGND VPWR VPWR U$$1792/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_667 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput90 b[32] VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__buf_6
XFILLER_123_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_72_2 dadda_fa_4_72_2/A dadda_fa_4_72_2/B dadda_fa_4_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_73_0/CIN dadda_fa_5_72_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_88_2 U$$2444/X U$$2577/X U$$2710/X VGND VGND VPWR VPWR dadda_fa_2_89_4/A
+ dadda_fa_2_88_5/B sky130_fd_sc_hd__fa_1
XFILLER_115_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_65_1 dadda_fa_4_65_1/A dadda_fa_4_65_1/B dadda_fa_4_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/B dadda_fa_5_65_1/B sky130_fd_sc_hd__fa_1
XFILLER_66_1076 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_42_0 dadda_fa_7_42_0/A dadda_fa_7_42_0/B dadda_fa_7_42_0/CIN VGND VGND
+ VPWR VPWR _339_/D _210_/D sky130_fd_sc_hd__fa_2
XFILLER_118_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_58_0 dadda_fa_4_58_0/A dadda_fa_4_58_0/B dadda_fa_4_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/A dadda_fa_5_58_1/A sky130_fd_sc_hd__fa_1
XTAP_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$410 final_adder.U$$414/B final_adder.U$$410/B VGND VGND VPWR VPWR
+ final_adder.U$$534/B sky130_fd_sc_hd__and2_1
XTAP_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$421 final_adder.U$$420/B final_adder.U$$299/X final_adder.U$$295/X
+ VGND VGND VPWR VPWR final_adder.U$$421/X sky130_fd_sc_hd__a21o_1
XTAP_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$432 final_adder.U$$436/B final_adder.U$$432/B VGND VGND VPWR VPWR
+ final_adder.U$$556/B sky130_fd_sc_hd__and2_1
XTAP_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$443 final_adder.U$$442/B final_adder.U$$321/X final_adder.U$$317/X
+ VGND VGND VPWR VPWR final_adder.U$$443/X sky130_fd_sc_hd__a21o_1
XTAP_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$454 final_adder.U$$458/B final_adder.U$$454/B VGND VGND VPWR VPWR
+ final_adder.U$$578/B sky130_fd_sc_hd__and2_1
XTAP_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$465 final_adder.U$$464/B final_adder.U$$343/X final_adder.U$$339/X
+ VGND VGND VPWR VPWR final_adder.U$$465/X sky130_fd_sc_hd__a21o_1
XU$$304 U$$578/A1 U$$316/A2 U$$717/A1 U$$316/B2 VGND VGND VPWR VPWR U$$305/A sky130_fd_sc_hd__a22o_1
XTAP_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$476 final_adder.U$$480/B final_adder.U$$476/B VGND VGND VPWR VPWR
+ final_adder.U$$600/B sky130_fd_sc_hd__and2_1
XTAP_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$315 U$$315/A U$$343/B VGND VGND VPWR VPWR U$$315/X sky130_fd_sc_hd__xor2_1
Xrepeater680 U$$527/B2 VGND VGND VPWR VPWR U$$473/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$487 final_adder.U$$486/B final_adder.U$$365/X final_adder.U$$361/X
+ VGND VGND VPWR VPWR final_adder.U$$487/X sky130_fd_sc_hd__a21o_1
XTAP_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$326 U$$461/B1 U$$350/A2 U$$54/A1 U$$350/B2 VGND VGND VPWR VPWR U$$327/A sky130_fd_sc_hd__a22o_1
Xrepeater691 U$$4238/B2 VGND VGND VPWR VPWR U$$4188/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$498 final_adder.U$$498/A final_adder.U$$498/B VGND VGND VPWR VPWR
+ final_adder.U$$614/A sky130_fd_sc_hd__and2_1
XTAP_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$337 U$$337/A U$$367/B VGND VGND VPWR VPWR U$$337/X sky130_fd_sc_hd__xor2_1
XU$$348 U$$483/B1 U$$350/A2 U$$76/A1 U$$350/B2 VGND VGND VPWR VPWR U$$349/A sky130_fd_sc_hd__a22o_1
XFILLER_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$359 U$$359/A U$$397/B VGND VGND VPWR VPWR U$$359/X sky130_fd_sc_hd__xor2_1
XFILLER_198_731 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_976 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1204 input65/X VGND VGND VPWR VPWR U$$4392/A1 sky130_fd_sc_hd__buf_6
XFILLER_154_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1215 U$$536/B VGND VGND VPWR VPWR U$$492/B sky130_fd_sc_hd__buf_6
XFILLER_181_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1226 U$$4382/B VGND VGND VPWR VPWR U$$4310/B sky130_fd_sc_hd__buf_6
Xrepeater1237 U$$4239/B VGND VGND VPWR VPWR U$$4189/B sky130_fd_sc_hd__buf_6
XFILLER_180_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1248 U$$410/A VGND VGND VPWR VPWR U$$395/B sky130_fd_sc_hd__buf_8
XFILLER_49_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1259 U$$3967/B VGND VGND VPWR VPWR U$$3947/B sky130_fd_sc_hd__buf_6
XFILLER_4_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_60_0 dadda_fa_3_60_0/A dadda_fa_3_60_0/B dadda_fa_3_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_0/B dadda_fa_4_60_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_76_0 dadda_fa_0_76_0/A U$$957/X U$$1090/X VGND VGND VPWR VPWR dadda_fa_1_77_8/B
+ dadda_fa_1_76_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$860 U$$860/A1 U$$892/A2 U$$860/B1 U$$892/B2 VGND VGND VPWR VPWR U$$861/A sky130_fd_sc_hd__a22o_1
XU$$1010 U$$1010/A U$$998/B VGND VGND VPWR VPWR U$$1010/X sky130_fd_sc_hd__xor2_1
XU$$871 U$$871/A U$$877/B VGND VGND VPWR VPWR U$$871/X sky130_fd_sc_hd__xor2_1
XU$$1021 U$$62/A1 U$$993/A2 U$$62/B1 U$$993/B2 VGND VGND VPWR VPWR U$$1022/A sky130_fd_sc_hd__a22o_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$882 U$$882/A1 U$$882/A2 U$$882/B1 U$$882/B2 VGND VGND VPWR VPWR U$$883/A sky130_fd_sc_hd__a22o_1
XU$$893 U$$893/A U$$929/B VGND VGND VPWR VPWR U$$893/X sky130_fd_sc_hd__xor2_1
XFILLER_56_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1032 U$$1032/A U$$1084/B VGND VGND VPWR VPWR U$$1032/X sky130_fd_sc_hd__xor2_1
XFILLER_90_386 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1043 U$$84/A1 U$$965/A2 U$$84/B1 U$$965/B2 VGND VGND VPWR VPWR U$$1044/A sky130_fd_sc_hd__a22o_1
XFILLER_32_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1054 U$$1054/A U$$1084/B VGND VGND VPWR VPWR U$$1054/X sky130_fd_sc_hd__xor2_1
XFILLER_177_915 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1065 U$$2709/A1 U$$963/X U$$2709/B1 U$$964/X VGND VGND VPWR VPWR U$$1066/A sky130_fd_sc_hd__a22o_1
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1076 U$$1076/A U$$1076/B VGND VGND VPWR VPWR U$$1076/X sky130_fd_sc_hd__xor2_1
XFILLER_204_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1087 U$$2318/B1 U$$1093/A2 U$$952/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1088/A
+ sky130_fd_sc_hd__a22o_1
XU$$1098 U$$1205/B VGND VGND VPWR VPWR U$$1098/Y sky130_fd_sc_hd__inv_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_82_1 dadda_fa_5_82_1/A dadda_fa_5_82_1/B dadda_fa_5_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_83_0/B dadda_fa_7_82_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_98_1 U$$2730/X U$$2863/X U$$2996/X VGND VGND VPWR VPWR dadda_fa_3_99_1/A
+ dadda_fa_3_98_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_75_0 dadda_fa_5_75_0/A dadda_fa_5_75_0/B dadda_fa_5_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_76_0/A dadda_fa_6_75_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_74_8 dadda_fa_1_74_8/A dadda_fa_1_74_8/B dadda_fa_1_74_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_75_3/A dadda_fa_3_74_0/A sky130_fd_sc_hd__fa_1
XFILLER_140_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_67_7 dadda_fa_1_67_7/A dadda_fa_1_67_7/B dadda_fa_1_67_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_2/CIN dadda_fa_2_67_5/CIN sky130_fd_sc_hd__fa_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_93_0 U$$2054/Y U$$2188/X U$$2321/X VGND VGND VPWR VPWR dadda_fa_2_94_5/A
+ dadda_fa_2_93_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3907 U$$3907/A U$$3909/B VGND VGND VPWR VPWR U$$3907/X sky130_fd_sc_hd__xor2_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$240 final_adder.U$$240/A final_adder.U$$240/B VGND VGND VPWR VPWR
+ final_adder.U$$368/B sky130_fd_sc_hd__and2_1
XTAP_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$251 final_adder.U$$5/SUM final_adder.U$$4/COUT final_adder.U$$5/COUT
+ VGND VGND VPWR VPWR final_adder.U$$251/X sky130_fd_sc_hd__a21o_1
XU$$3918 U$$4466/A1 U$$3926/A2 U$$4466/B1 U$$3926/B2 VGND VGND VPWR VPWR U$$3919/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3929 U$$3929/A U$$3947/B VGND VGND VPWR VPWR U$$3929/X sky130_fd_sc_hd__xor2_1
XTAP_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$101 U$$101/A U$$111/B VGND VGND VPWR VPWR U$$101/X sky130_fd_sc_hd__xor2_1
XFILLER_100_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$262 final_adder.U$$264/B final_adder.U$$262/B VGND VGND VPWR VPWR
+ final_adder.U$$388/B sky130_fd_sc_hd__and2_1
Xdadda_fa_6_105_0 dadda_fa_6_105_0/A dadda_fa_6_105_0/B dadda_fa_6_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_106_0/B dadda_fa_7_105_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$273 final_adder.U$$272/B final_adder.U$$147/X final_adder.U$$145/X
+ VGND VGND VPWR VPWR final_adder.U$$273/X sky130_fd_sc_hd__a21o_1
XTAP_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$112 U$$384/B1 U$$122/A2 U$$251/A1 U$$122/B2 VGND VGND VPWR VPWR U$$113/A sky130_fd_sc_hd__a22o_1
XTAP_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$284 final_adder.U$$286/B final_adder.U$$284/B VGND VGND VPWR VPWR
+ final_adder.U$$410/B sky130_fd_sc_hd__and2_1
XTAP_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$123 U$$123/A U$$127/B VGND VGND VPWR VPWR U$$123/X sky130_fd_sc_hd__xor2_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$295 final_adder.U$$294/B final_adder.U$$169/X final_adder.U$$167/X
+ VGND VGND VPWR VPWR final_adder.U$$295/X sky130_fd_sc_hd__a21o_1
XTAP_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$134 U$$817/B1 U$$134/A2 U$$134/B1 U$$134/B2 VGND VGND VPWR VPWR U$$135/A sky130_fd_sc_hd__a22o_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$145 U$$8/A1 U$$165/A2 U$$8/B1 U$$165/B2 VGND VGND VPWR VPWR U$$146/A sky130_fd_sc_hd__a22o_1
XFILLER_150_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$156 U$$156/A U$$160/B VGND VGND VPWR VPWR U$$156/X sky130_fd_sc_hd__xor2_1
XTAP_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_25_3 dadda_fa_3_25_3/A dadda_fa_3_25_3/B dadda_fa_3_25_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_26_1/B dadda_fa_4_25_2/CIN sky130_fd_sc_hd__fa_1
XU$$167 U$$578/A1 U$$175/A2 U$$32/A1 U$$175/B2 VGND VGND VPWR VPWR U$$168/A sky130_fd_sc_hd__a22o_1
XTAP_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$178 U$$178/A U$$184/B VGND VGND VPWR VPWR U$$178/X sky130_fd_sc_hd__xor2_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$189 U$$598/B1 U$$217/A2 U$$54/A1 U$$217/B2 VGND VGND VPWR VPWR U$$190/A sky130_fd_sc_hd__a22o_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_550 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_395_ _399_/CLK _395_/D VGND VGND VPWR VPWR _395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_92_0 dadda_fa_6_92_0/A dadda_fa_6_92_0/B dadda_fa_6_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_93_0/B dadda_fa_7_92_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_138_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1001 U$$2123/A1 VGND VGND VPWR VPWR U$$342/A1 sky130_fd_sc_hd__buf_4
Xrepeater1012 U$$3300/A1 VGND VGND VPWR VPWR U$$3026/A1 sky130_fd_sc_hd__buf_4
XFILLER_153_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1023 input86/X VGND VGND VPWR VPWR U$$4311/B1 sky130_fd_sc_hd__buf_6
Xrepeater1034 U$$2391/A1 VGND VGND VPWR VPWR U$$62/A1 sky130_fd_sc_hd__buf_4
Xrepeater1045 U$$3485/A1 VGND VGND VPWR VPWR U$$3483/B1 sky130_fd_sc_hd__buf_6
Xrepeater1056 input82/X VGND VGND VPWR VPWR U$$4442/A1 sky130_fd_sc_hd__buf_6
Xrepeater1067 input80/X VGND VGND VPWR VPWR U$$3614/B1 sky130_fd_sc_hd__buf_8
Xrepeater1078 U$$4297/B1 VGND VGND VPWR VPWR U$$461/B1 sky130_fd_sc_hd__buf_4
XFILLER_107_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1089 input78/X VGND VGND VPWR VPWR U$$50/A1 sky130_fd_sc_hd__buf_6
XFILLER_141_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_124_0_1870 VGND VGND VPWR VPWR dadda_fa_5_124_0/A dadda_fa_5_124_0_1870/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_96_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1040 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$690 U$$688/B U$$685/A input2/X U$$685/Y VGND VGND VPWR VPWR U$$690/X sky130_fd_sc_hd__a22o_4
XFILLER_211_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1091 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_222 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_80_8 U$$4290/X U$$4423/X VGND VGND VPWR VPWR dadda_fa_2_81_3/B dadda_fa_3_80_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1590 U$$2717/A1 VGND VGND VPWR VPWR U$$2032/A1 sky130_fd_sc_hd__buf_4
XFILLER_8_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_72_5 U$$4008/X U$$4141/X U$$4274/X VGND VGND VPWR VPWR dadda_fa_2_73_2/A
+ dadda_fa_2_72_5/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_65_4 U$$4127/X U$$4260/X U$$4393/X VGND VGND VPWR VPWR dadda_fa_2_66_1/CIN
+ dadda_fa_2_65_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_3 U$$2783/X U$$2916/X U$$3049/X VGND VGND VPWR VPWR dadda_fa_2_59_1/B
+ dadda_fa_2_58_4/B sky130_fd_sc_hd__fa_1
XFILLER_67_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_35_2 dadda_fa_4_35_2/A dadda_fa_4_35_2/B dadda_fa_4_35_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_36_0/CIN dadda_fa_5_35_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_28_1 dadda_fa_4_28_1/A dadda_fa_4_28_1/B dadda_fa_4_28_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/B dadda_fa_5_28_1/B sky130_fd_sc_hd__fa_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_180_ _314_/CLK _180_/D VGND VGND VPWR VPWR _180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4405 U$$4405/A U$$4405/B VGND VGND VPWR VPWR U$$4405/X sky130_fd_sc_hd__xor2_1
XFILLER_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4416 input68/X U$$4388/X input69/X U$$4498/B2 VGND VGND VPWR VPWR U$$4417/A sky130_fd_sc_hd__a22o_1
XTAP_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_60_3 U$$1324/X U$$1457/X U$$1590/X VGND VGND VPWR VPWR dadda_fa_1_61_7/A
+ dadda_fa_1_60_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4427 U$$4427/A U$$4427/B VGND VGND VPWR VPWR U$$4427/X sky130_fd_sc_hd__xor2_1
XU$$4438 U$$4438/A1 U$$4388/X U$$4440/A1 U$$4389/X VGND VGND VPWR VPWR U$$4439/A sky130_fd_sc_hd__a22o_1
XFILLER_65_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_3_17_1 U$$440/X U$$573/X VGND VGND VPWR VPWR dadda_fa_4_18_1/CIN dadda_ha_3_17_1/SUM
+ sky130_fd_sc_hd__ha_1
XU$$4449 U$$4449/A U$$4449/B VGND VGND VPWR VPWR U$$4449/X sky130_fd_sc_hd__xor2_1
XU$$3704 U$$3702/B input49/X input50/X U$$3699/Y VGND VGND VPWR VPWR U$$3704/X sky130_fd_sc_hd__a22o_2
XTAP_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3715 U$$3852/A1 U$$3753/A2 U$$3852/B1 U$$3753/B2 VGND VGND VPWR VPWR U$$3716/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3726 U$$3726/A U$$3740/B VGND VGND VPWR VPWR U$$3726/X sky130_fd_sc_hd__xor2_1
XTAP_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_73 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_448 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3737 U$$3737/A1 U$$3739/A2 U$$3737/B1 U$$3739/B2 VGND VGND VPWR VPWR U$$3738/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_30_1 input180/X dadda_fa_3_30_1/B dadda_fa_3_30_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_31_0/CIN dadda_fa_4_30_2/A sky130_fd_sc_hd__fa_1
XU$$3748 U$$3748/A U$$3754/B VGND VGND VPWR VPWR U$$3748/X sky130_fd_sc_hd__xor2_1
XTAP_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3759 input83/X U$$3703/X U$$3761/A1 U$$3777/B2 VGND VGND VPWR VPWR U$$3760/A sky130_fd_sc_hd__a22o_1
XTAP_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_23_0 U$$319/X U$$452/X U$$585/X VGND VGND VPWR VPWR dadda_fa_4_24_0/B
+ dadda_fa_4_23_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_378_ _384_/CLK _378_/D VGND VGND VPWR VPWR _378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_82_4 dadda_fa_2_82_4/A dadda_fa_2_82_4/B dadda_fa_2_82_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_1/CIN dadda_fa_3_82_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_138_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_75_3 dadda_fa_2_75_3/A dadda_fa_2_75_3/B dadda_fa_2_75_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/B dadda_fa_3_75_3/B sky130_fd_sc_hd__fa_1
Xdadda_fa_2_68_2 dadda_fa_2_68_2/A dadda_fa_2_68_2/B dadda_fa_2_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/A dadda_fa_3_68_3/A sky130_fd_sc_hd__fa_1
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_45_1 dadda_fa_5_45_1/A dadda_fa_5_45_1/B dadda_fa_5_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_46_0/B dadda_fa_7_45_0/A sky130_fd_sc_hd__fa_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_38_0 dadda_fa_5_38_0/A dadda_fa_5_38_0/B dadda_fa_5_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_39_0/A dadda_fa_6_38_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_504 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_112_0 dadda_fa_5_112_0/A dadda_fa_5_112_0/B dadda_fa_5_112_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_113_0/A dadda_fa_6_112_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_30_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_1151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_70_2 U$$3073/X U$$3206/X U$$3339/X VGND VGND VPWR VPWR dadda_fa_2_71_1/A
+ dadda_fa_2_70_4/A sky130_fd_sc_hd__fa_1
XFILLER_115_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_1 U$$2793/X U$$2926/X U$$3059/X VGND VGND VPWR VPWR dadda_fa_2_64_0/CIN
+ dadda_fa_2_63_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_927 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_40_0 dadda_fa_4_40_0/A dadda_fa_4_40_0/B dadda_fa_4_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/A dadda_fa_5_40_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_1_56_0 U$$1183/X U$$1316/X U$$1449/X VGND VGND VPWR VPWR dadda_fa_2_57_0/B
+ dadda_fa_2_56_3/B sky130_fd_sc_hd__fa_1
XFILLER_75_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_971 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1609 U$$2292/B1 U$$1637/A2 U$$2568/B1 U$$1637/B2 VGND VGND VPWR VPWR U$$1610/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_610 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_301_ _304_/CLK _301_/D VGND VGND VPWR VPWR _301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$408_1759 VGND VGND VPWR VPWR U$$408_1759/HI U$$408/B1 sky130_fd_sc_hd__conb_1
XFILLER_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_232_ _362_/CLK _232_/D VGND VGND VPWR VPWR _232_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_92_3 dadda_fa_3_92_3/A dadda_fa_3_92_3/B dadda_fa_3_92_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_93_1/B dadda_fa_4_92_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_136_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_85_2 dadda_fa_3_85_2/A dadda_fa_3_85_2/B dadda_fa_3_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_1/A dadda_fa_4_85_2/B sky130_fd_sc_hd__fa_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_78_1 dadda_fa_3_78_1/A dadda_fa_3_78_1/B dadda_fa_3_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_0/CIN dadda_fa_4_78_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_55_0 dadda_fa_6_55_0/A dadda_fa_6_55_0/B dadda_fa_6_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_56_0/B dadda_fa_7_55_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater509 U$$3118/A2 VGND VGND VPWR VPWR U$$3082/A2 sky130_fd_sc_hd__buf_12
XFILLER_78_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4202 input101/X U$$4226/A2 input102/X U$$4226/B2 VGND VGND VPWR VPWR U$$4203/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4213 U$$4213/A U$$4227/B VGND VGND VPWR VPWR U$$4213/X sky130_fd_sc_hd__xor2_1
XU$$4224 input113/X U$$4240/A2 U$$4500/A1 U$$4240/B2 VGND VGND VPWR VPWR U$$4225/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4235 U$$4235/A U$$4239/B VGND VGND VPWR VPWR U$$4235/X sky130_fd_sc_hd__xor2_1
XFILLER_66_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3501 U$$3775/A1 U$$3503/A2 U$$3775/B1 U$$3503/B2 VGND VGND VPWR VPWR U$$3502/A
+ sky130_fd_sc_hd__a22o_1
XU$$4246 U$$4246/A VGND VGND VPWR VPWR U$$4246/Y sky130_fd_sc_hd__inv_1
XU$$4257 U$$4394/A1 U$$4275/A2 U$$4396/A1 U$$4275/B2 VGND VGND VPWR VPWR U$$4258/A
+ sky130_fd_sc_hd__a22o_1
XU$$3512 U$$3512/A U$$3518/B VGND VGND VPWR VPWR U$$3512/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_114_2 dadda_fa_4_114_2/A dadda_fa_4_114_2/B dadda_ha_3_114_1/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_115_0/CIN dadda_fa_5_114_1/CIN sky130_fd_sc_hd__fa_1
XU$$3523 U$$783/A1 U$$3527/A2 U$$783/B1 U$$3527/B2 VGND VGND VPWR VPWR U$$3524/A sky130_fd_sc_hd__a22o_1
XFILLER_1_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4268 U$$4268/A U$$4310/B VGND VGND VPWR VPWR U$$4268/X sky130_fd_sc_hd__xor2_1
XU$$3534 U$$3534/A U$$3550/B VGND VGND VPWR VPWR U$$3534/X sky130_fd_sc_hd__xor2_1
XU$$4279 input68/X U$$4327/A2 U$$32/B1 U$$4327/B2 VGND VGND VPWR VPWR U$$4280/A sky130_fd_sc_hd__a22o_1
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3545 U$$3545/A1 U$$3549/A2 U$$3684/A1 U$$3549/B2 VGND VGND VPWR VPWR U$$3546/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2800 U$$4442/B1 U$$2844/A2 U$$3211/B1 U$$2844/B2 VGND VGND VPWR VPWR U$$2801/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2811 U$$2811/A U$$2817/B VGND VGND VPWR VPWR U$$2811/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_107_1 dadda_fa_4_107_1/A dadda_fa_4_107_1/B dadda_fa_4_107_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/B dadda_fa_5_107_1/B sky130_fd_sc_hd__fa_1
XU$$3556 U$$3556/A U$$3561/A VGND VGND VPWR VPWR U$$3556/X sky130_fd_sc_hd__xor2_1
XFILLER_34_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2822 input95/X U$$2858/A2 U$$3646/A1 U$$2858/B2 VGND VGND VPWR VPWR U$$2823/A
+ sky130_fd_sc_hd__a22o_1
XU$$3567 U$$3565/B input47/X input48/X U$$3562/Y VGND VGND VPWR VPWR U$$3567/X sky130_fd_sc_hd__a22o_4
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3578 U$$3578/A1 U$$3612/A2 U$$3578/B1 U$$3612/B2 VGND VGND VPWR VPWR U$$3579/A
+ sky130_fd_sc_hd__a22o_1
XU$$2833 U$$2833/A U$$2837/B VGND VGND VPWR VPWR U$$2833/X sky130_fd_sc_hd__xor2_1
XFILLER_92_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3589 U$$3589/A U$$3613/B VGND VGND VPWR VPWR U$$3589/X sky130_fd_sc_hd__xor2_1
XU$$2844 U$$3116/B1 U$$2844/A2 U$$2981/B1 U$$2844/B2 VGND VGND VPWR VPWR U$$2845/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2855 U$$2855/A U$$2859/B VGND VGND VPWR VPWR U$$2855/X sky130_fd_sc_hd__xor2_1
XFILLER_61_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2866 U$$3414/A1 U$$2868/A2 U$$3414/B1 U$$2868/B2 VGND VGND VPWR VPWR U$$2867/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_160 U$$2957/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2877 input36/X VGND VGND VPWR VPWR U$$2877/Y sky130_fd_sc_hd__inv_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2888 U$$2888/A U$$2922/B VGND VGND VPWR VPWR U$$2888/X sky130_fd_sc_hd__xor2_1
XFILLER_33_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_171 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2899 U$$981/A1 U$$2919/A2 U$$709/A1 U$$2919/B2 VGND VGND VPWR VPWR U$$2900/A sky130_fd_sc_hd__a22o_1
XANTENNA_193 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_80_1 dadda_fa_2_80_1/A dadda_fa_2_80_1/B dadda_fa_2_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_0/CIN dadda_fa_3_80_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_73_0 dadda_fa_2_73_0/A dadda_fa_2_73_0/B dadda_fa_2_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_0/B dadda_fa_3_73_2/B sky130_fd_sc_hd__fa_1
XFILLER_114_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$817 final_adder.U$$784/A final_adder.U$$737/X final_adder.U$$705/X
+ VGND VGND VPWR VPWR final_adder.U$$817/X sky130_fd_sc_hd__a21o_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4449_1801 VGND VGND VPWR VPWR U$$4449_1801/HI U$$4449/B sky130_fd_sc_hd__conb_1
XFILLER_57_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$839 final_adder.U$$742/X final_adder.U$$807/X final_adder.U$$743/X
+ VGND VGND VPWR VPWR final_adder.U$$839/X sky130_fd_sc_hd__a21o_2
XFILLER_151_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_79 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_95_1 dadda_fa_4_95_1/A dadda_fa_4_95_1/B dadda_fa_4_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/B dadda_fa_5_95_1/B sky130_fd_sc_hd__fa_1
XFILLER_119_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_72_0 dadda_fa_7_72_0/A dadda_fa_7_72_0/B dadda_fa_7_72_0/CIN VGND VGND
+ VPWR VPWR _369_/D _240_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_88_0 dadda_fa_4_88_0/A dadda_fa_4_88_0/B dadda_fa_4_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/A dadda_fa_5_88_1/A sky130_fd_sc_hd__fa_1
XFILLER_180_559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_109_3 U$$4348/X U$$4481/X input139/X VGND VGND VPWR VPWR dadda_fa_4_110_1/B
+ dadda_fa_4_109_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput370 output370/A VGND VGND VPWR VPWR o[87] sky130_fd_sc_hd__buf_2
Xoutput381 output381/A VGND VGND VPWR VPWR o[97] sky130_fd_sc_hd__buf_2
XFILLER_156_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4389_1770 VGND VGND VPWR VPWR U$$4389_1770/HI U$$4389/B1 sky130_fd_sc_hd__conb_1
XFILLER_210_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2107 U$$3749/B1 U$$2113/A2 U$$3614/B1 U$$2113/B2 VGND VGND VPWR VPWR U$$2108/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_727 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2118 U$$2118/A U$$2150/B VGND VGND VPWR VPWR U$$2118/X sky130_fd_sc_hd__xor2_1
XU$$2129 U$$896/A1 U$$2169/A2 U$$896/B1 U$$2169/B2 VGND VGND VPWR VPWR U$$2130/A sky130_fd_sc_hd__a22o_1
XFILLER_28_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1023 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1406 U$$719/B1 U$$1448/A2 U$$312/A1 U$$1448/B2 VGND VGND VPWR VPWR U$$1407/A sky130_fd_sc_hd__a22o_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1417 U$$1417/A U$$1423/B VGND VGND VPWR VPWR U$$1417/X sky130_fd_sc_hd__xor2_1
XFILLER_167_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1428 U$$56/B1 U$$1434/A2 U$$2661/B1 U$$1434/B2 VGND VGND VPWR VPWR U$$1429/A sky130_fd_sc_hd__a22o_1
XU$$1439 U$$1439/A U$$1449/B VGND VGND VPWR VPWR U$$1439/X sky130_fd_sc_hd__xor2_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_215_ _218_/CLK _215_/D VGND VGND VPWR VPWR _215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_90_0 dadda_fa_3_90_0/A dadda_fa_3_90_0/B dadda_fa_3_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_0/B dadda_fa_4_90_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_137_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_52_5 dadda_fa_2_52_5/A dadda_fa_2_52_5/B dadda_fa_2_52_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_53_2/A dadda_fa_4_52_0/A sky130_fd_sc_hd__fa_2
XU$$4010 U$$4010/A U$$4044/B VGND VGND VPWR VPWR U$$4010/X sky130_fd_sc_hd__xor2_1
XFILLER_65_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4021 input77/X U$$4107/A2 input78/X U$$4107/B2 VGND VGND VPWR VPWR U$$4022/A sky130_fd_sc_hd__a22o_1
XFILLER_211_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4032 U$$4032/A U$$4036/B VGND VGND VPWR VPWR U$$4032/X sky130_fd_sc_hd__xor2_1
XU$$4043 U$$4043/A1 U$$4043/A2 U$$4043/B1 U$$4043/B2 VGND VGND VPWR VPWR U$$4044/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4054 U$$4054/A U$$4080/B VGND VGND VPWR VPWR U$$4054/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_45_4 dadda_fa_2_45_4/A dadda_fa_2_45_4/B dadda_fa_2_45_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_1/CIN dadda_fa_3_45_3/CIN sky130_fd_sc_hd__fa_1
XU$$3320 U$$4005/A1 U$$3320/A2 U$$4144/A1 U$$3320/B2 VGND VGND VPWR VPWR U$$3321/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4065 U$$4476/A1 U$$4077/A2 U$$4476/B1 U$$4077/B2 VGND VGND VPWR VPWR U$$4066/A
+ sky130_fd_sc_hd__a22o_1
XU$$4076 U$$4076/A U$$4078/B VGND VGND VPWR VPWR U$$4076/X sky130_fd_sc_hd__xor2_1
XU$$3331 U$$3331/A U$$3375/B VGND VGND VPWR VPWR U$$3331/X sky130_fd_sc_hd__xor2_1
XFILLER_19_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4087 input113/X U$$4101/A2 U$$4361/B1 U$$4101/B2 VGND VGND VPWR VPWR U$$4088/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3342 U$$4027/A1 U$$3378/A2 U$$3344/A1 U$$3346/B2 VGND VGND VPWR VPWR U$$3343/A
+ sky130_fd_sc_hd__a22o_1
XU$$4098 U$$4098/A U$$4110/A VGND VGND VPWR VPWR U$$4098/X sky130_fd_sc_hd__xor2_1
XFILLER_19_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3353 U$$3353/A U$$3389/B VGND VGND VPWR VPWR U$$3353/X sky130_fd_sc_hd__xor2_1
XU$$3364 U$$3775/A1 U$$3292/X U$$3775/B1 U$$3293/X VGND VGND VPWR VPWR U$$3365/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_38_3 U$$2344/X U$$2477/X U$$2610/X VGND VGND VPWR VPWR dadda_fa_3_39_1/B
+ dadda_fa_3_38_3/B sky130_fd_sc_hd__fa_1
XFILLER_94_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2630 U$$2630/A U$$2658/B VGND VGND VPWR VPWR U$$2630/X sky130_fd_sc_hd__xor2_1
XFILLER_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3375 U$$3375/A U$$3375/B VGND VGND VPWR VPWR U$$3375/X sky130_fd_sc_hd__xor2_1
XU$$3386 U$$783/A1 U$$3388/A2 U$$783/B1 U$$3390/B2 VGND VGND VPWR VPWR U$$3387/A sky130_fd_sc_hd__a22o_1
XU$$2641 U$$312/A1 U$$2727/A2 U$$38/B1 U$$2727/B2 VGND VGND VPWR VPWR U$$2642/A sky130_fd_sc_hd__a22o_1
XU$$3397 U$$3397/A U$$3417/B VGND VGND VPWR VPWR U$$3397/X sky130_fd_sc_hd__xor2_1
XU$$2652 U$$2652/A U$$2658/B VGND VGND VPWR VPWR U$$2652/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2663 U$$3485/A1 U$$2691/A2 U$$3211/B1 U$$2691/B2 VGND VGND VPWR VPWR U$$2664/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2674 U$$2674/A U$$2680/B VGND VGND VPWR VPWR U$$2674/X sky130_fd_sc_hd__xor2_1
XU$$2685 U$$4055/A1 U$$2735/A2 U$$4055/B1 U$$2735/B2 VGND VGND VPWR VPWR U$$2686/A
+ sky130_fd_sc_hd__a22o_1
XU$$1940 U$$3447/A1 U$$1990/A2 U$$3584/B1 U$$1990/B2 VGND VGND VPWR VPWR U$$1941/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1951 U$$1951/A U$$1993/B VGND VGND VPWR VPWR U$$1951/X sky130_fd_sc_hd__xor2_1
XFILLER_61_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_906 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2696 U$$2696/A U$$2716/B VGND VGND VPWR VPWR U$$2696/X sky130_fd_sc_hd__xor2_1
XU$$1962 U$$3878/B1 U$$1990/A2 U$$731/A1 U$$1990/B2 VGND VGND VPWR VPWR U$$1963/A
+ sky130_fd_sc_hd__a22o_1
XU$$1973 U$$1973/A U$$2017/B VGND VGND VPWR VPWR U$$1973/X sky130_fd_sc_hd__xor2_1
XU$$1984 U$$1984/A1 U$$2016/A2 U$$2123/A1 U$$2016/B2 VGND VGND VPWR VPWR U$$1985/A
+ sky130_fd_sc_hd__a22o_1
XU$$4479_1816 VGND VGND VPWR VPWR U$$4479_1816/HI U$$4479/B sky130_fd_sc_hd__conb_1
XFILLER_166_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1995 U$$1995/A U$$2043/B VGND VGND VPWR VPWR U$$1995/X sky130_fd_sc_hd__xor2_1
XFILLER_193_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput109 b[4] VGND VGND VPWR VPWR input109/X sky130_fd_sc_hd__buf_8
XTAP_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$603 final_adder.U$$602/B final_adder.U$$487/X final_adder.U$$479/X
+ VGND VGND VPWR VPWR final_adder.U$$603/X sky130_fd_sc_hd__a21o_1
XTAP_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$614 final_adder.U$$614/A final_adder.U$$614/B VGND VGND VPWR VPWR
+ final_adder.U$$718/A sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$625 final_adder.U$$616/A final_adder.U$$255/X final_adder.U$$501/X
+ VGND VGND VPWR VPWR final_adder.U$$625/X sky130_fd_sc_hd__a21o_2
XFILLER_9_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$636 final_adder.U$$652/B final_adder.U$$636/B VGND VGND VPWR VPWR
+ final_adder.U$$748/B sky130_fd_sc_hd__and2_1
XTAP_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater840 U$$1649/X VGND VGND VPWR VPWR U$$1736/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$647 final_adder.U$$646/B final_adder.U$$543/X final_adder.U$$527/X
+ VGND VGND VPWR VPWR final_adder.U$$647/X sky130_fd_sc_hd__a21o_1
XTAP_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater851 U$$1591/B2 VGND VGND VPWR VPWR U$$1557/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$658 final_adder.U$$674/B final_adder.U$$658/B VGND VGND VPWR VPWR
+ final_adder.U$$770/B sky130_fd_sc_hd__and2_1
XTAP_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater862 U$$142/X VGND VGND VPWR VPWR U$$231/B2 sky130_fd_sc_hd__buf_6
XFILLER_84_554 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$669 final_adder.U$$668/B final_adder.U$$565/X final_adder.U$$549/X
+ VGND VGND VPWR VPWR final_adder.U$$669/X sky130_fd_sc_hd__a21o_1
XU$$508 U$$508/A U$$528/B VGND VGND VPWR VPWR U$$508/X sky130_fd_sc_hd__xor2_1
Xrepeater873 U$$1238/X VGND VGND VPWR VPWR U$$1367/B2 sky130_fd_sc_hd__buf_4
Xrepeater884 U$$1101/X VGND VGND VPWR VPWR U$$1230/B2 sky130_fd_sc_hd__buf_6
XU$$519 U$$654/B1 U$$521/A2 U$$521/A1 U$$521/B2 VGND VGND VPWR VPWR U$$520/A sky130_fd_sc_hd__a22o_1
XFILLER_38_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater895 U$$4430/B2 VGND VGND VPWR VPWR U$$4426/B2 sky130_fd_sc_hd__buf_6
XFILLER_38_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$80 U$$80/A1 U$$80/A2 U$$82/A1 U$$80/B2 VGND VGND VPWR VPWR U$$81/A sky130_fd_sc_hd__a22o_1
XU$$91 U$$91/A U$$99/B VGND VGND VPWR VPWR U$$91/X sky130_fd_sc_hd__xor2_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_60 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_82 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_93 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1408 U$$2170/B VGND VGND VPWR VPWR U$$2150/B sky130_fd_sc_hd__buf_6
XFILLER_115_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1419 input22/X VGND VGND VPWR VPWR U$$2047/B sky130_fd_sc_hd__buf_6
XFILLER_197_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_107_0 U$$3413/X U$$3546/X U$$3679/X VGND VGND VPWR VPWR dadda_fa_4_108_0/B
+ dadda_fa_4_107_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_55_3 dadda_fa_3_55_3/A dadda_fa_3_55_3/B dadda_fa_3_55_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_56_1/B dadda_fa_4_55_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_48_2 dadda_fa_3_48_2/A dadda_fa_3_48_2/B dadda_fa_3_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_1/A dadda_fa_4_48_2/B sky130_fd_sc_hd__fa_1
XFILLER_101_191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_18_0 dadda_fa_6_18_0/A dadda_fa_6_18_0/B dadda_fa_6_18_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_19_0/B dadda_fa_7_18_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_16_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1203 U$$1203/A U$$1205/B VGND VGND VPWR VPWR U$$1203/X sky130_fd_sc_hd__xor2_1
XFILLER_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1214 U$$527/B1 U$$1230/A2 U$$2449/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1215/A
+ sky130_fd_sc_hd__a22o_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1225 U$$1225/A U$$1232/A VGND VGND VPWR VPWR U$$1225/X sky130_fd_sc_hd__xor2_1
XFILLER_204_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1236 U$$1338/B U$$1236/B VGND VGND VPWR VPWR U$$1236/X sky130_fd_sc_hd__and2_1
XFILLER_16_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1247 U$$2069/A1 U$$1271/A2 U$$2206/B1 U$$1271/B2 VGND VGND VPWR VPWR U$$1248/A
+ sky130_fd_sc_hd__a22o_1
XU$$1258 U$$1258/A U$$1270/B VGND VGND VPWR VPWR U$$1258/X sky130_fd_sc_hd__xor2_1
XU$$1269 U$$719/B1 U$$1271/A2 U$$721/B1 U$$1271/B2 VGND VGND VPWR VPWR U$$1270/A sky130_fd_sc_hd__a22o_1
XFILLER_203_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1030 final_adder.U$$6/SUM final_adder.U$$505/X VGND VGND VPWR VPWR
+ output351/A sky130_fd_sc_hd__xor2_1
XFILLER_8_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1041 final_adder.U$$238/B final_adder.U$$1041/B VGND VGND VPWR VPWR
+ output293/A sky130_fd_sc_hd__xor2_1
XFILLER_184_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1052 final_adder.U$$226/A final_adder.U$$727/X VGND VGND VPWR VPWR
+ output305/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1063 final_adder.U$$216/B final_adder.U$$987/X VGND VGND VPWR VPWR
+ output317/A sky130_fd_sc_hd__xor2_1
XFILLER_176_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1074 final_adder.U$$204/A final_adder.U$$817/X VGND VGND VPWR VPWR
+ output330/A sky130_fd_sc_hd__xor2_1
XFILLER_176_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1085 final_adder.U$$194/B final_adder.U$$965/X VGND VGND VPWR VPWR
+ output342/A sky130_fd_sc_hd__xor2_1
XFILLER_171_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1096 final_adder.U$$182/A final_adder.U$$891/X VGND VGND VPWR VPWR
+ output354/A sky130_fd_sc_hd__xor2_1
XFILLER_171_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_50_2 dadda_fa_2_50_2/A dadda_fa_2_50_2/B dadda_fa_2_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/A dadda_fa_3_50_3/A sky130_fd_sc_hd__fa_1
XFILLER_61_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_43_1 U$$2354/X U$$2487/X U$$2620/X VGND VGND VPWR VPWR dadda_fa_3_44_0/CIN
+ dadda_fa_3_43_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_20_0 dadda_fa_5_20_0/A dadda_fa_5_20_0/B dadda_fa_5_20_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_21_0/A dadda_fa_6_20_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3150 U$$3150/A VGND VGND VPWR VPWR U$$3150/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_2_36_0 U$$744/X U$$877/X U$$1010/X VGND VGND VPWR VPWR dadda_fa_3_37_0/B
+ dadda_fa_3_36_2/B sky130_fd_sc_hd__fa_1
XFILLER_4_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3161 U$$3296/B1 U$$3187/A2 U$$3300/A1 U$$3187/B2 VGND VGND VPWR VPWR U$$3162/A
+ sky130_fd_sc_hd__a22o_1
XU$$3172 U$$3172/A U$$3264/B VGND VGND VPWR VPWR U$$3172/X sky130_fd_sc_hd__xor2_1
XFILLER_81_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3183 U$$3183/A1 U$$3187/A2 U$$3183/B1 U$$3187/B2 VGND VGND VPWR VPWR U$$3184/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3194 U$$3194/A U$$3208/B VGND VGND VPWR VPWR U$$3194/X sky130_fd_sc_hd__xor2_1
XU$$2460 U$$2460/A U$$2465/A VGND VGND VPWR VPWR U$$2460/X sky130_fd_sc_hd__xor2_1
XU$$2471 U$$2469/B U$$2466/A input30/X U$$2466/Y VGND VGND VPWR VPWR U$$2471/X sky130_fd_sc_hd__a22o_4
XFILLER_59_1084 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2482 U$$2754/B1 U$$2490/A2 U$$2621/A1 U$$2490/B2 VGND VGND VPWR VPWR U$$2483/A
+ sky130_fd_sc_hd__a22o_1
XU$$2493 U$$2493/A U$$2525/B VGND VGND VPWR VPWR U$$2493/X sky130_fd_sc_hd__xor2_1
XFILLER_195_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1770 U$$948/A1 U$$1770/A2 U$$2044/B1 U$$1770/B2 VGND VGND VPWR VPWR U$$1771/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1781 input18/X VGND VGND VPWR VPWR U$$1781/Y sky130_fd_sc_hd__inv_1
XFILLER_107_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1792 U$$1792/A U$$1820/B VGND VGND VPWR VPWR U$$1792/X sky130_fd_sc_hd__xor2_1
XFILLER_194_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_537 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput80 b[23] VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__buf_12
XFILLER_174_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput91 b[33] VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__buf_8
XFILLER_122_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_23 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_88_3 U$$2843/X U$$2976/X U$$3109/X VGND VGND VPWR VPWR dadda_fa_2_89_4/B
+ dadda_fa_2_88_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_157_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_65_2 dadda_fa_4_65_2/A dadda_fa_4_65_2/B dadda_fa_4_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_66_0/CIN dadda_fa_5_65_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_58_1 dadda_fa_4_58_1/A dadda_fa_4_58_1/B dadda_fa_4_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/B dadda_fa_5_58_1/B sky130_fd_sc_hd__fa_1
XTAP_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$400 final_adder.U$$404/B final_adder.U$$400/B VGND VGND VPWR VPWR
+ final_adder.U$$524/B sky130_fd_sc_hd__and2_1
XFILLER_190_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$411 final_adder.U$$410/B final_adder.U$$289/X final_adder.U$$285/X
+ VGND VGND VPWR VPWR final_adder.U$$411/X sky130_fd_sc_hd__a21o_1
XTAP_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_35_0 dadda_fa_7_35_0/A dadda_fa_7_35_0/B dadda_fa_7_35_0/CIN VGND VGND
+ VPWR VPWR _332_/D _203_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$422 final_adder.U$$426/B final_adder.U$$422/B VGND VGND VPWR VPWR
+ final_adder.U$$546/B sky130_fd_sc_hd__and2_1
XTAP_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$433 final_adder.U$$432/B final_adder.U$$311/X final_adder.U$$307/X
+ VGND VGND VPWR VPWR final_adder.U$$433/X sky130_fd_sc_hd__a21o_1
XTAP_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$444 final_adder.U$$448/B final_adder.U$$444/B VGND VGND VPWR VPWR
+ final_adder.U$$568/B sky130_fd_sc_hd__and2_1
XTAP_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$455 final_adder.U$$454/B final_adder.U$$333/X final_adder.U$$329/X
+ VGND VGND VPWR VPWR final_adder.U$$455/X sky130_fd_sc_hd__a21o_1
XTAP_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$466 final_adder.U$$470/B final_adder.U$$466/B VGND VGND VPWR VPWR
+ final_adder.U$$590/B sky130_fd_sc_hd__and2_1
XU$$305 U$$305/A U$$379/B VGND VGND VPWR VPWR U$$305/X sky130_fd_sc_hd__xor2_1
XTAP_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater670 U$$4297/B2 VGND VGND VPWR VPWR U$$4275/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$477 final_adder.U$$476/B final_adder.U$$355/X final_adder.U$$351/X
+ VGND VGND VPWR VPWR final_adder.U$$477/X sky130_fd_sc_hd__a21o_1
Xrepeater681 U$$515/B2 VGND VGND VPWR VPWR U$$437/B2 sky130_fd_sc_hd__buf_4
XTAP_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$316 U$$42/A1 U$$316/A2 U$$44/A1 U$$316/B2 VGND VGND VPWR VPWR U$$317/A sky130_fd_sc_hd__a22o_1
XFILLER_57_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$488 final_adder.U$$492/B final_adder.U$$488/B VGND VGND VPWR VPWR
+ final_adder.U$$612/B sky130_fd_sc_hd__and2_1
XTAP_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$327 U$$327/A U$$351/B VGND VGND VPWR VPWR U$$327/X sky130_fd_sc_hd__xor2_1
Xrepeater692 U$$4240/B2 VGND VGND VPWR VPWR U$$4238/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$499 final_adder.U$$498/B final_adder.U$$377/X final_adder.U$$373/X
+ VGND VGND VPWR VPWR final_adder.U$$499/X sky130_fd_sc_hd__a21o_1
XU$$338 U$$610/B1 U$$366/A2 U$$66/A1 U$$366/B2 VGND VGND VPWR VPWR U$$339/A sky130_fd_sc_hd__a22o_1
XU$$349 U$$349/A U$$351/B VGND VGND VPWR VPWR U$$349/X sky130_fd_sc_hd__xor2_1
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1048 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1205 U$$637/B VGND VGND VPWR VPWR U$$607/B sky130_fd_sc_hd__buf_6
XFILLER_148_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1216 U$$546/B VGND VGND VPWR VPWR U$$536/B sky130_fd_sc_hd__buf_4
XFILLER_5_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1227 U$$4370/B VGND VGND VPWR VPWR U$$4330/B sky130_fd_sc_hd__buf_6
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1238 U$$4247/A VGND VGND VPWR VPWR U$$4239/B sky130_fd_sc_hd__buf_6
Xrepeater1249 U$$410/A VGND VGND VPWR VPWR U$$411/A sky130_fd_sc_hd__buf_4
XFILLER_180_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_60_1 dadda_fa_3_60_1/A dadda_fa_3_60_1/B dadda_fa_3_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_0/CIN dadda_fa_4_60_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_53_0 dadda_fa_3_53_0/A dadda_fa_3_53_0/B dadda_fa_3_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_0/B dadda_fa_4_53_1/CIN sky130_fd_sc_hd__fa_2
XFILLER_0_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_69_0 U$$410/Y U$$544/X U$$677/X VGND VGND VPWR VPWR dadda_fa_1_70_6/A
+ dadda_fa_1_69_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$850 U$$850/A1 U$$872/A2 U$$850/B1 U$$872/B2 VGND VGND VPWR VPWR U$$851/A sky130_fd_sc_hd__a22o_1
XFILLER_169_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$861 U$$861/A U$$929/B VGND VGND VPWR VPWR U$$861/X sky130_fd_sc_hd__xor2_1
XU$$1000 U$$999/X U$$996/B VGND VGND VPWR VPWR U$$1000/X sky130_fd_sc_hd__xor2_1
XU$$1011 U$$598/B1 U$$997/A2 U$$54/A1 U$$997/B2 VGND VGND VPWR VPWR U$$1012/A sky130_fd_sc_hd__a22o_1
XFILLER_90_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$872 U$$48/B1 U$$872/A2 U$$52/A1 U$$872/B2 VGND VGND VPWR VPWR U$$873/A sky130_fd_sc_hd__a22o_1
XU$$1022 U$$1022/A U$$994/B VGND VGND VPWR VPWR U$$1022/X sky130_fd_sc_hd__xor2_1
XU$$883 U$$883/A U$$883/B VGND VGND VPWR VPWR U$$883/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$894 U$$894/A1 U$$938/A2 U$$896/A1 U$$938/B2 VGND VGND VPWR VPWR U$$895/A sky130_fd_sc_hd__a22o_1
XFILLER_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1033 U$$483/B1 U$$1057/A2 U$$76/A1 U$$1057/B2 VGND VGND VPWR VPWR U$$1034/A sky130_fd_sc_hd__a22o_1
XFILLER_204_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1044 U$$1044/A U$$968/B VGND VGND VPWR VPWR U$$1044/X sky130_fd_sc_hd__xor2_1
XFILLER_50_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_398 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1055 U$$96/A1 U$$1057/A2 U$$98/A1 U$$1057/B2 VGND VGND VPWR VPWR U$$1056/A sky130_fd_sc_hd__a22o_1
XFILLER_188_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1066 U$$1066/A U$$962/A VGND VGND VPWR VPWR U$$1066/X sky130_fd_sc_hd__xor2_1
XFILLER_177_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1077 U$$527/B1 U$$1083/A2 U$$942/A1 U$$1083/B2 VGND VGND VPWR VPWR U$$1078/A sky130_fd_sc_hd__a22o_1
XU$$1088 U$$1088/A U$$1095/A VGND VGND VPWR VPWR U$$1088/X sky130_fd_sc_hd__xor2_1
XU$$1099 U$$1209/B U$$1099/B VGND VGND VPWR VPWR U$$1099/X sky130_fd_sc_hd__and2_1
XFILLER_143_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_110_0 dadda_fa_7_110_0/A dadda_fa_7_110_0/B dadda_fa_7_110_0/CIN VGND
+ VGND VPWR VPWR _407_/D _278_/D sky130_fd_sc_hd__fa_1
XFILLER_185_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_98_2 U$$3129/X U$$3262/X U$$3395/X VGND VGND VPWR VPWR dadda_fa_3_99_1/B
+ dadda_fa_3_98_3/A sky130_fd_sc_hd__fa_1
XFILLER_172_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_75_1 dadda_fa_5_75_1/A dadda_fa_5_75_1/B dadda_fa_5_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_76_0/B dadda_fa_7_75_0/A sky130_fd_sc_hd__fa_1
XFILLER_104_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_68_0 dadda_fa_5_68_0/A dadda_fa_5_68_0/B dadda_fa_5_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_69_0/A dadda_fa_6_68_0/CIN sky130_fd_sc_hd__fa_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_67_8 dadda_fa_1_67_8/A dadda_fa_1_67_8/B dadda_fa_1_67_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_68_3/A dadda_fa_3_67_0/A sky130_fd_sc_hd__fa_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_310 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_7_0 dadda_fa_6_7_0/A dadda_fa_6_7_0/B dadda_fa_6_7_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_8_0/B dadda_fa_7_7_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_179_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2290 U$$4480/B1 U$$2326/A2 U$$3114/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2291/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_297 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1002 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_93_1 U$$2454/X U$$2587/X U$$2720/X VGND VGND VPWR VPWR dadda_fa_2_94_5/B
+ dadda_fa_3_93_0/A sky130_fd_sc_hd__fa_1
XFILLER_190_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_70_0 dadda_fa_4_70_0/A dadda_fa_4_70_0/B dadda_fa_4_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/A dadda_fa_5_70_1/A sky130_fd_sc_hd__fa_1
XFILLER_1_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_86_0 dadda_fa_1_86_0/A U$$1642/X U$$1775/X VGND VGND VPWR VPWR dadda_fa_2_87_2/CIN
+ dadda_fa_2_86_4/B sky130_fd_sc_hd__fa_1
XFILLER_150_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_2_106_1 U$$3278/X U$$3411/X VGND VGND VPWR VPWR dadda_fa_3_107_3/CIN dadda_fa_4_106_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$230 final_adder.U$$230/A final_adder.U$$230/B VGND VGND VPWR VPWR
+ final_adder.U$$358/B sky130_fd_sc_hd__and2_1
XFILLER_182_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3908 U$$4043/B1 U$$3840/X U$$3908/B1 U$$3841/X VGND VGND VPWR VPWR U$$3909/A sky130_fd_sc_hd__a22o_1
XFILLER_92_619 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$241 final_adder.U$$240/B final_adder.U$$241/A2 final_adder.U$$241/B1
+ VGND VGND VPWR VPWR final_adder.U$$241/X sky130_fd_sc_hd__a21o_1
XTAP_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3919 U$$3919/A U$$3927/B VGND VGND VPWR VPWR U$$3919/X sky130_fd_sc_hd__xor2_1
XTAP_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$252 final_adder.U$$252/A final_adder.U$$3/SUM VGND VGND VPWR VPWR
+ final_adder.U$$378/A sky130_fd_sc_hd__and2_1
XTAP_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$263 final_adder.U$$262/B final_adder.U$$137/X final_adder.U$$135/X
+ VGND VGND VPWR VPWR final_adder.U$$263/X sky130_fd_sc_hd__a21o_1
XTAP_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$102 U$$787/A1 U$$134/A2 U$$926/A1 U$$134/B2 VGND VGND VPWR VPWR U$$103/A sky130_fd_sc_hd__a22o_1
XFILLER_100_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$274 final_adder.U$$276/B final_adder.U$$274/B VGND VGND VPWR VPWR
+ final_adder.U$$400/B sky130_fd_sc_hd__and2_1
XU$$113 U$$113/A U$$127/B VGND VGND VPWR VPWR U$$113/X sky130_fd_sc_hd__xor2_1
XTAP_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$285 final_adder.U$$284/B final_adder.U$$159/X final_adder.U$$157/X
+ VGND VGND VPWR VPWR final_adder.U$$285/X sky130_fd_sc_hd__a21o_1
XFILLER_205_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$124 U$$944/B1 U$$134/A2 U$$811/A1 U$$134/B2 VGND VGND VPWR VPWR U$$125/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$296 final_adder.U$$298/B final_adder.U$$296/B VGND VGND VPWR VPWR
+ final_adder.U$$422/B sky130_fd_sc_hd__and2_1
XTAP_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$135 U$$135/A U$$3/A VGND VGND VPWR VPWR U$$135/X sky130_fd_sc_hd__xor2_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$146 U$$146/A U$$160/B VGND VGND VPWR VPWR U$$146/X sky130_fd_sc_hd__xor2_1
XTAP_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$157 U$$20/A1 U$$165/A2 U$$22/A1 U$$165/B2 VGND VGND VPWR VPWR U$$158/A sky130_fd_sc_hd__a22o_1
XTAP_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$168 U$$168/A U$$184/B VGND VGND VPWR VPWR U$$168/X sky130_fd_sc_hd__xor2_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$179 U$$179/A1 U$$209/A2 U$$866/A1 U$$209/B2 VGND VGND VPWR VPWR U$$180/A sky130_fd_sc_hd__a22o_1
XFILLER_150_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_394_ _394_/CLK _394_/D VGND VGND VPWR VPWR _394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_85_0 dadda_fa_6_85_0/A dadda_fa_6_85_0/B dadda_fa_6_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_86_0/B dadda_fa_7_85_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1002 U$$4452/A1 VGND VGND VPWR VPWR U$$2123/A1 sky130_fd_sc_hd__buf_6
Xrepeater1013 input87/X VGND VGND VPWR VPWR U$$4396/A1 sky130_fd_sc_hd__buf_4
Xrepeater1024 U$$610/B1 VGND VGND VPWR VPWR U$$64/A1 sky130_fd_sc_hd__buf_4
XFILLER_175_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1035 U$$610/A1 VGND VGND VPWR VPWR U$$2391/A1 sky130_fd_sc_hd__buf_4
XFILLER_154_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1046 U$$4442/B1 VGND VGND VPWR VPWR U$$4307/A1 sky130_fd_sc_hd__buf_6
Xrepeater1057 U$$741/A1 VGND VGND VPWR VPWR U$$56/A1 sky130_fd_sc_hd__buf_4
Xrepeater1068 U$$874/B1 VGND VGND VPWR VPWR U$$328/A1 sky130_fd_sc_hd__buf_4
Xrepeater1079 U$$4297/B1 VGND VGND VPWR VPWR U$$4436/A1 sky130_fd_sc_hd__buf_6
XFILLER_141_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1020 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$680 U$$954/A1 U$$552/X U$$956/A1 U$$553/X VGND VGND VPWR VPWR U$$681/A sky130_fd_sc_hd__a22o_1
XU$$691 U$$691/A1 U$$711/A2 U$$967/A1 U$$711/B2 VGND VGND VPWR VPWR U$$692/A sky130_fd_sc_hd__a22o_1
XFILLER_147_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1239_1713 VGND VGND VPWR VPWR U$$1239_1713/HI U$$1239/A1 sky130_fd_sc_hd__conb_1
XFILLER_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1580 input114/X VGND VGND VPWR VPWR U$$116/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_67_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1591 U$$4498/A1 VGND VGND VPWR VPWR U$$2717/A1 sky130_fd_sc_hd__buf_4
XFILLER_8_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1036 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_72_6 U$$4407/X input226/X dadda_fa_1_72_6/CIN VGND VGND VPWR VPWR dadda_fa_2_73_2/B
+ dadda_fa_2_72_5/B sky130_fd_sc_hd__fa_1
XFILLER_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_65_5 input218/X dadda_fa_1_65_5/B dadda_fa_1_65_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_66_2/A dadda_fa_2_65_5/A sky130_fd_sc_hd__fa_1
XFILLER_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_58_4 U$$3182/X U$$3315/X U$$3448/X VGND VGND VPWR VPWR dadda_fa_2_59_1/CIN
+ dadda_fa_2_58_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_28_2 dadda_fa_4_28_2/A dadda_fa_4_28_2/B dadda_fa_4_28_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_29_0/CIN dadda_fa_5_28_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4406 U$$4406/A1 U$$4388/X U$$4408/A1 U$$4430/B2 VGND VGND VPWR VPWR U$$4407/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4417 U$$4417/A U$$4417/B VGND VGND VPWR VPWR U$$4417/X sky130_fd_sc_hd__xor2_1
XFILLER_93_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4428 U$$4428/A1 U$$4388/X U$$4430/A1 U$$4430/B2 VGND VGND VPWR VPWR U$$4429/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4439 U$$4439/A U$$4439/B VGND VGND VPWR VPWR U$$4439/X sky130_fd_sc_hd__xor2_1
XFILLER_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3705 U$$3705/A1 U$$3793/A2 U$$3979/B1 U$$3793/B2 VGND VGND VPWR VPWR U$$3706/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3716 U$$3716/A U$$3754/B VGND VGND VPWR VPWR U$$3716/X sky130_fd_sc_hd__xor2_1
XTAP_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3727 U$$4275/A1 U$$3739/A2 U$$3727/B1 U$$3739/B2 VGND VGND VPWR VPWR U$$3728/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3738 U$$3738/A U$$3774/B VGND VGND VPWR VPWR U$$3738/X sky130_fd_sc_hd__xor2_1
XFILLER_206_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3749 U$$3749/A1 U$$3793/A2 U$$3749/B1 U$$3793/B2 VGND VGND VPWR VPWR U$$3750/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1778_1722 VGND VGND VPWR VPWR U$$1778_1722/HI U$$1778/B1 sky130_fd_sc_hd__conb_1
XFILLER_45_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_30_2 dadda_fa_3_30_2/A dadda_fa_3_30_2/B dadda_fa_3_30_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_31_1/A dadda_fa_4_30_2/B sky130_fd_sc_hd__fa_1
XFILLER_205_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_23_1 U$$718/X U$$851/X U$$984/X VGND VGND VPWR VPWR dadda_fa_4_24_0/CIN
+ dadda_fa_4_23_2/A sky130_fd_sc_hd__fa_1
XFILLER_73_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_16_0 U$$39/X U$$172/X U$$305/X VGND VGND VPWR VPWR dadda_fa_4_17_1/CIN
+ dadda_fa_4_16_2/B sky130_fd_sc_hd__fa_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_377_ _377_/CLK _377_/D VGND VGND VPWR VPWR _377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_82_5 dadda_fa_2_82_5/A dadda_fa_2_82_5/B dadda_fa_2_82_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_83_2/A dadda_fa_4_82_0/A sky130_fd_sc_hd__fa_2
XFILLER_126_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_75_4 dadda_fa_2_75_4/A dadda_fa_2_75_4/B dadda_fa_2_75_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_1/CIN dadda_fa_3_75_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_68_3 dadda_fa_2_68_3/A dadda_fa_2_68_3/B dadda_fa_2_68_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/B dadda_fa_3_68_3/B sky130_fd_sc_hd__fa_1
XFILLER_68_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_38_1 dadda_fa_5_38_1/A dadda_fa_5_38_1/B dadda_fa_5_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_39_0/B dadda_fa_7_38_0/A sky130_fd_sc_hd__fa_2
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_112_1 dadda_fa_5_112_1/A dadda_fa_5_112_1/B dadda_fa_5_112_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_113_0/B dadda_fa_7_112_0/A sky130_fd_sc_hd__fa_1
XFILLER_166_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_105_0 dadda_fa_5_105_0/A dadda_fa_5_105_0/B dadda_fa_5_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_106_0/A dadda_fa_6_105_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_70_3 U$$3472/X U$$3605/X U$$3738/X VGND VGND VPWR VPWR dadda_fa_2_71_1/B
+ dadda_fa_2_70_4/B sky130_fd_sc_hd__fa_1
XFILLER_113_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_2 U$$3192/X U$$3325/X U$$3458/X VGND VGND VPWR VPWR dadda_fa_2_64_1/A
+ dadda_fa_2_63_4/A sky130_fd_sc_hd__fa_1
XFILLER_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_40_1 dadda_fa_4_40_1/A dadda_fa_4_40_1/B dadda_fa_4_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/B dadda_fa_5_40_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_56_1 U$$1582/X U$$1715/X U$$1848/X VGND VGND VPWR VPWR dadda_fa_2_57_0/CIN
+ dadda_fa_2_56_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_33_0 dadda_fa_4_33_0/A dadda_fa_4_33_0/B dadda_fa_4_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/A dadda_fa_5_33_1/A sky130_fd_sc_hd__fa_1
XFILLER_28_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_49_0 U$$105/X U$$238/X U$$371/X VGND VGND VPWR VPWR dadda_fa_2_50_0/CIN
+ dadda_fa_2_49_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_41_1197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_983 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_300_ _304_/CLK _300_/D VGND VGND VPWR VPWR _300_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_231_ _360_/CLK _231_/D VGND VGND VPWR VPWR _231_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_85_3 dadda_fa_3_85_3/A dadda_fa_3_85_3/B dadda_fa_3_85_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_86_1/B dadda_fa_4_85_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_156_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_78_2 dadda_fa_3_78_2/A dadda_fa_3_78_2/B dadda_fa_3_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_1/A dadda_fa_4_78_2/B sky130_fd_sc_hd__fa_1
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_48_0 dadda_fa_6_48_0/A dadda_fa_6_48_0/B dadda_fa_6_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_49_0/B dadda_fa_7_48_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_120_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4203 U$$4203/A U$$4227/B VGND VGND VPWR VPWR U$$4203/X sky130_fd_sc_hd__xor2_1
XFILLER_133_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4214 U$$4488/A1 U$$4226/A2 U$$4490/A1 U$$4226/B2 VGND VGND VPWR VPWR U$$4215/A
+ sky130_fd_sc_hd__a22o_1
XU$$4225 U$$4225/A U$$4247/A VGND VGND VPWR VPWR U$$4225/X sky130_fd_sc_hd__xor2_1
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4236 U$$4236/A1 U$$4238/A2 U$$4512/A1 U$$4238/B2 VGND VGND VPWR VPWR U$$4237/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3502 U$$3502/A U$$3504/B VGND VGND VPWR VPWR U$$3502/X sky130_fd_sc_hd__xor2_1
XU$$4247 U$$4247/A VGND VGND VPWR VPWR U$$4247/Y sky130_fd_sc_hd__inv_1
XU$$3513 U$$3648/B1 U$$3517/A2 U$$4335/B1 U$$3517/B2 VGND VGND VPWR VPWR U$$3514/A
+ sky130_fd_sc_hd__a22o_1
XU$$4258 U$$4258/A U$$4278/B VGND VGND VPWR VPWR U$$4258/X sky130_fd_sc_hd__xor2_1
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3524 U$$3524/A U$$3528/B VGND VGND VPWR VPWR U$$3524/X sky130_fd_sc_hd__xor2_1
XU$$4269 U$$4269/A1 U$$4275/A2 U$$4269/B1 U$$4275/B2 VGND VGND VPWR VPWR U$$4270/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3535 input111/X U$$3559/A2 input112/X U$$3559/B2 VGND VGND VPWR VPWR U$$3536/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3546 U$$3546/A U$$3550/B VGND VGND VPWR VPWR U$$3546/X sky130_fd_sc_hd__xor2_1
XU$$2801 U$$2801/A U$$2837/B VGND VGND VPWR VPWR U$$2801/X sky130_fd_sc_hd__xor2_1
XU$$3557 U$$4103/B1 U$$3559/A2 U$$3557/B1 U$$3559/B2 VGND VGND VPWR VPWR U$$3558/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2812 U$$4045/A1 U$$2828/A2 U$$3088/A1 U$$2828/B2 VGND VGND VPWR VPWR U$$2813/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_107_2 dadda_fa_4_107_2/A dadda_fa_4_107_2/B dadda_fa_4_107_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_108_0/CIN dadda_fa_5_107_1/CIN sky130_fd_sc_hd__fa_1
XU$$2823 U$$2823/A U$$2859/B VGND VGND VPWR VPWR U$$2823/X sky130_fd_sc_hd__xor2_1
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3568 U$$3568/A1 U$$3612/A2 U$$3979/B1 U$$3612/B2 VGND VGND VPWR VPWR U$$3569/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2834 U$$2834/A1 U$$2844/A2 U$$3108/B1 U$$2844/B2 VGND VGND VPWR VPWR U$$2835/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3579 U$$3579/A U$$3609/B VGND VGND VPWR VPWR U$$3579/X sky130_fd_sc_hd__xor2_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2845 U$$2845/A U$$2845/B VGND VGND VPWR VPWR U$$2845/X sky130_fd_sc_hd__xor2_1
XFILLER_206_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2856 U$$388/B1 U$$2868/A2 U$$3680/A1 U$$2868/B2 VGND VGND VPWR VPWR U$$2857/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_110 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2867 U$$2867/A U$$2869/B VGND VGND VPWR VPWR U$$2867/X sky130_fd_sc_hd__xor2_1
XANTENNA_150 U$$3227/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_161 U$$2810/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2878 input37/X VGND VGND VPWR VPWR U$$2880/B sky130_fd_sc_hd__inv_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2889 U$$3026/A1 U$$2921/A2 U$$3028/A1 U$$2921/B2 VGND VGND VPWR VPWR U$$2890/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_502 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_80_2 dadda_fa_2_80_2/A dadda_fa_2_80_2/B dadda_fa_2_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/A dadda_fa_3_80_3/A sky130_fd_sc_hd__fa_1
XFILLER_142_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_73_1 dadda_fa_2_73_1/A dadda_fa_2_73_1/B dadda_fa_2_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_0/CIN dadda_fa_3_73_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_50_0 dadda_fa_5_50_0/A dadda_fa_5_50_0/B dadda_fa_5_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_51_0/A dadda_fa_6_50_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_66_0 dadda_fa_2_66_0/A dadda_fa_2_66_0/B dadda_fa_2_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_0/B dadda_fa_3_66_2/B sky130_fd_sc_hd__fa_1
XFILLER_69_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$807 final_adder.U$$774/A final_adder.U$$727/X final_adder.U$$695/X
+ VGND VGND VPWR VPWR final_adder.U$$807/X sky130_fd_sc_hd__a21o_1
XFILLER_151_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$829 final_adder.U$$796/A final_adder.U$$505/X final_adder.U$$717/X
+ VGND VGND VPWR VPWR final_adder.U$$829/X sky130_fd_sc_hd__a21o_1
XFILLER_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 a[0] VGND VGND VPWR VPWR U$$1/A sky130_fd_sc_hd__buf_2
XFILLER_99_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_clk _239_/CLK VGND VGND VPWR VPWR _368_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4421_1787 VGND VGND VPWR VPWR U$$4421_1787/HI U$$4421/B sky130_fd_sc_hd__conb_1
Xdadda_fa_4_95_2 dadda_fa_4_95_2/A dadda_fa_4_95_2/B dadda_fa_4_95_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_96_0/CIN dadda_fa_5_95_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_153_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_974 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_88_1 dadda_fa_4_88_1/A dadda_fa_4_88_1/B dadda_fa_4_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/B dadda_fa_5_88_1/B sky130_fd_sc_hd__fa_1
XFILLER_161_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_65_0 dadda_fa_7_65_0/A dadda_fa_7_65_0/B dadda_fa_7_65_0/CIN VGND VGND
+ VPWR VPWR _362_/D _233_/D sky130_fd_sc_hd__fa_1
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput360 output360/A VGND VGND VPWR VPWR o[78] sky130_fd_sc_hd__buf_2
XFILLER_0_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput371 output371/A VGND VGND VPWR VPWR o[88] sky130_fd_sc_hd__buf_2
Xoutput382 output382/A VGND VGND VPWR VPWR o[98] sky130_fd_sc_hd__buf_2
XFILLER_126_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_39_clk _239_/CLK VGND VGND VPWR VPWR _379_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$2108 U$$2108/A U$$2114/B VGND VGND VPWR VPWR U$$2108/X sky130_fd_sc_hd__xor2_1
XU$$2119 U$$3213/B1 U$$2149/A2 U$$477/A1 U$$2149/B2 VGND VGND VPWR VPWR U$$2120/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1407 U$$1407/A U$$1449/B VGND VGND VPWR VPWR U$$1407/X sky130_fd_sc_hd__xor2_1
XU$$1418 U$$594/B1 U$$1470/A2 U$$461/A1 U$$1470/B2 VGND VGND VPWR VPWR U$$1419/A sky130_fd_sc_hd__a22o_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1429 U$$1429/A U$$1459/B VGND VGND VPWR VPWR U$$1429/X sky130_fd_sc_hd__xor2_1
XFILLER_71_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_214_ _219_/CLK _214_/D VGND VGND VPWR VPWR _214_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_11_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_90_1 dadda_fa_3_90_1/A dadda_fa_3_90_1/B dadda_fa_3_90_1/CIN VGND VGND
+ VPWR VPWR ANTENNA_0/DIODE dadda_fa_4_90_2/A sky130_fd_sc_hd__fa_2
XFILLER_13_1085 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_83_0 dadda_fa_3_83_0/A dadda_fa_3_83_0/B dadda_fa_3_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_0/B dadda_fa_4_83_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4000 U$$4000/A U$$4036/B VGND VGND VPWR VPWR U$$4000/X sky130_fd_sc_hd__xor2_1
XFILLER_120_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4011 U$$4011/A1 U$$4011/A2 U$$4011/B1 U$$4011/B2 VGND VGND VPWR VPWR U$$4012/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4022 U$$4022/A input55/X VGND VGND VPWR VPWR U$$4022/X sky130_fd_sc_hd__xor2_1
XFILLER_120_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4033 U$$4307/A1 U$$4035/A2 U$$4309/A1 U$$4035/B2 VGND VGND VPWR VPWR U$$4034/A
+ sky130_fd_sc_hd__a22o_1
XU$$4044 U$$4044/A U$$4044/B VGND VGND VPWR VPWR U$$4044/X sky130_fd_sc_hd__xor2_1
XU$$3310 input126/X U$$3394/A2 input127/X U$$3394/B2 VGND VGND VPWR VPWR U$$3311/A
+ sky130_fd_sc_hd__a22o_1
XU$$4055 U$$4055/A1 U$$4079/A2 U$$4055/B1 U$$4079/B2 VGND VGND VPWR VPWR U$$4056/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_1170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4066 U$$4066/A U$$4078/B VGND VGND VPWR VPWR U$$4066/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_0 U$$4354/X U$$4487/X input143/X VGND VGND VPWR VPWR dadda_fa_5_113_0/A
+ dadda_fa_5_112_1/A sky130_fd_sc_hd__fa_1
XFILLER_20_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_45_5 dadda_fa_2_45_5/A dadda_fa_2_45_5/B dadda_fa_2_45_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_46_2/A dadda_fa_4_45_0/A sky130_fd_sc_hd__fa_1
XFILLER_47_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3321 U$$3321/A U$$3321/B VGND VGND VPWR VPWR U$$3321/X sky130_fd_sc_hd__xor2_1
XU$$4077 U$$4488/A1 U$$4077/A2 U$$4077/B1 U$$4077/B2 VGND VGND VPWR VPWR U$$4078/A
+ sky130_fd_sc_hd__a22o_1
XU$$3332 U$$4428/A1 U$$3374/A2 U$$4430/A1 U$$3374/B2 VGND VGND VPWR VPWR U$$3333/A
+ sky130_fd_sc_hd__a22o_1
XU$$3343 U$$3343/A U$$3425/A VGND VGND VPWR VPWR U$$3343/X sky130_fd_sc_hd__xor2_1
XFILLER_93_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4088 U$$4088/A U$$4110/A VGND VGND VPWR VPWR U$$4088/X sky130_fd_sc_hd__xor2_1
XU$$4099 U$$4236/A1 U$$4103/A2 U$$4099/B1 U$$4103/B2 VGND VGND VPWR VPWR U$$4100/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_38_4 U$$2624/B input188/X dadda_fa_2_38_4/CIN VGND VGND VPWR VPWR dadda_fa_3_39_1/CIN
+ dadda_fa_3_38_3/CIN sky130_fd_sc_hd__fa_1
XU$$3354 U$$4311/B1 U$$3388/A2 U$$3356/A1 U$$3390/B2 VGND VGND VPWR VPWR U$$3355/A
+ sky130_fd_sc_hd__a22o_1
XU$$2620 U$$2620/A U$$2624/B VGND VGND VPWR VPWR U$$2620/X sky130_fd_sc_hd__xor2_1
XU$$3365 U$$3365/A U$$3377/B VGND VGND VPWR VPWR U$$3365/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3376 U$$3376/A1 U$$3292/X U$$3378/A1 U$$3293/X VGND VGND VPWR VPWR U$$3377/A sky130_fd_sc_hd__a22o_1
XU$$2631 U$$711/B1 U$$2653/A2 U$$578/A1 U$$2653/B2 VGND VGND VPWR VPWR U$$2632/A sky130_fd_sc_hd__a22o_1
XU$$2642 U$$2642/A U$$2650/B VGND VGND VPWR VPWR U$$2642/X sky130_fd_sc_hd__xor2_1
XU$$3387 U$$3387/A U$$3389/B VGND VGND VPWR VPWR U$$3387/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2653 U$$3884/B1 U$$2653/A2 U$$3612/B1 U$$2653/B2 VGND VGND VPWR VPWR U$$2654/A
+ sky130_fd_sc_hd__a22o_1
XU$$3398 U$$3944/B1 U$$3416/A2 U$$384/B1 U$$3416/B2 VGND VGND VPWR VPWR U$$3399/A
+ sky130_fd_sc_hd__a22o_1
XU$$2664 U$$2664/A U$$2680/B VGND VGND VPWR VPWR U$$2664/X sky130_fd_sc_hd__xor2_1
XU$$2675 U$$2810/B1 U$$2683/A2 U$$3088/A1 U$$2683/B2 VGND VGND VPWR VPWR U$$2676/A
+ sky130_fd_sc_hd__a22o_1
XU$$1930 U$$2065/B1 U$$1990/A2 U$$2343/A1 U$$1990/B2 VGND VGND VPWR VPWR U$$1931/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2686 U$$2686/A U$$2739/A VGND VGND VPWR VPWR U$$2686/X sky130_fd_sc_hd__xor2_1
XU$$1941 U$$1941/A U$$1991/B VGND VGND VPWR VPWR U$$1941/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1952 U$$993/A1 U$$1960/A2 U$$993/B1 U$$1960/B2 VGND VGND VPWR VPWR U$$1953/A sky130_fd_sc_hd__a22o_1
XU$$2697 U$$3245/A1 U$$2711/A2 U$$3245/B1 U$$2711/B2 VGND VGND VPWR VPWR U$$2698/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1963 U$$1963/A U$$1991/B VGND VGND VPWR VPWR U$$1963/X sky130_fd_sc_hd__xor2_1
XFILLER_210_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1974 U$$3481/A1 U$$2016/A2 U$$3618/B1 U$$2016/B2 VGND VGND VPWR VPWR U$$1975/A
+ sky130_fd_sc_hd__a22o_1
XU$$1985 U$$1985/A U$$2017/B VGND VGND VPWR VPWR U$$1985/X sky130_fd_sc_hd__xor2_1
XU$$1996 U$$3366/A1 U$$2040/A2 U$$3366/B1 U$$2040/B2 VGND VGND VPWR VPWR U$$1997/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_98_0 dadda_fa_5_98_0/A dadda_fa_5_98_0/B dadda_fa_5_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_99_0/A dadda_fa_6_98_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_147_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$604 final_adder.U$$612/B final_adder.U$$604/B VGND VGND VPWR VPWR
+ final_adder.U$$708/A sky130_fd_sc_hd__and2_1
XFILLER_96_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$615 final_adder.U$$614/B final_adder.U$$499/X final_adder.U$$491/X
+ VGND VGND VPWR VPWR final_adder.U$$615/X sky130_fd_sc_hd__a21o_1
XFILLER_116_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater830 U$$1923/X VGND VGND VPWR VPWR U$$2046/B2 sky130_fd_sc_hd__buf_6
XFILLER_56_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$637 final_adder.U$$636/B final_adder.U$$533/X final_adder.U$$517/X
+ VGND VGND VPWR VPWR final_adder.U$$637/X sky130_fd_sc_hd__a21o_1
XTAP_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater841 U$$1746/B2 VGND VGND VPWR VPWR U$$1696/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$648 final_adder.U$$664/B final_adder.U$$648/B VGND VGND VPWR VPWR
+ final_adder.U$$760/B sky130_fd_sc_hd__and2_1
XTAP_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater852 U$$1607/B2 VGND VGND VPWR VPWR U$$1591/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$659 final_adder.U$$658/B final_adder.U$$555/X final_adder.U$$539/X
+ VGND VGND VPWR VPWR final_adder.U$$659/X sky130_fd_sc_hd__a21o_1
XFILLER_45_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater863 U$$1502/B2 VGND VGND VPWR VPWR U$$1448/B2 sky130_fd_sc_hd__buf_4
XFILLER_56_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$509 U$$920/A1 U$$521/A2 U$$783/B1 U$$521/B2 VGND VGND VPWR VPWR U$$510/A sky130_fd_sc_hd__a22o_1
Xrepeater874 U$$1238/X VGND VGND VPWR VPWR U$$1349/B2 sky130_fd_sc_hd__buf_6
XFILLER_84_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater885 U$$1204/B2 VGND VGND VPWR VPWR U$$1162/B2 sky130_fd_sc_hd__buf_4
Xrepeater896 U$$4432/B2 VGND VGND VPWR VPWR U$$4430/B2 sky130_fd_sc_hd__buf_6
XFILLER_72_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$70 U$$70/A1 U$$80/A2 U$$72/A1 U$$80/B2 VGND VGND VPWR VPWR U$$71/A sky130_fd_sc_hd__a22o_1
XFILLER_53_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$81 U$$81/A U$$81/B VGND VGND VPWR VPWR U$$81/X sky130_fd_sc_hd__xor2_1
XFILLER_198_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$92 U$$92/A1 U$$94/A2 U$$94/A1 U$$94/B2 VGND VGND VPWR VPWR U$$93/A sky130_fd_sc_hd__a22o_1
XFILLER_73_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_50 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_61 _342_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_72 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_83 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_94 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1409 U$$2178/B VGND VGND VPWR VPWR U$$2170/B sky130_fd_sc_hd__buf_12
XFILLER_181_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_107_1 U$$3812/X U$$3945/X U$$4078/X VGND VGND VPWR VPWR dadda_fa_4_108_0/CIN
+ dadda_fa_4_107_2/A sky130_fd_sc_hd__fa_1
XFILLER_180_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_48_3 dadda_fa_3_48_3/A dadda_fa_3_48_3/B dadda_fa_3_48_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_49_1/B dadda_fa_4_48_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_972 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1204 U$$2709/B1 U$$1204/A2 U$$932/A1 U$$1204/B2 VGND VGND VPWR VPWR U$$1205/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1215 U$$1215/A U$$1232/A VGND VGND VPWR VPWR U$$1215/X sky130_fd_sc_hd__xor2_1
XFILLER_188_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1226 U$$952/A1 U$$1230/A2 U$$2324/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1227/A
+ sky130_fd_sc_hd__a22o_1
XU$$1237 U$$1235/Y input10/X input9/X U$$1236/X U$$1233/Y VGND VGND VPWR VPWR U$$1237/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_71_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1248 U$$1248/A U$$1272/B VGND VGND VPWR VPWR U$$1248/X sky130_fd_sc_hd__xor2_1
XFILLER_188_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1259 U$$985/A1 U$$1289/A2 U$$2220/A1 U$$1291/B2 VGND VGND VPWR VPWR U$$1260/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1031 final_adder.U$$7/SUM final_adder.U$$1031/B VGND VGND VPWR VPWR
+ output362/A sky130_fd_sc_hd__xor2_1
XFILLER_156_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1042 final_adder.U$$236/A final_adder.U$$737/X VGND VGND VPWR VPWR
+ output294/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1053 final_adder.U$$226/B final_adder.U$$997/X VGND VGND VPWR VPWR
+ output306/A sky130_fd_sc_hd__xor2_1
XFILLER_184_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1064 final_adder.U$$214/A final_adder.U$$827/X VGND VGND VPWR VPWR
+ output319/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1075 final_adder.U$$204/B final_adder.U$$975/X VGND VGND VPWR VPWR
+ output331/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1086 final_adder.U$$192/A final_adder.U$$805/X VGND VGND VPWR VPWR
+ output343/A sky130_fd_sc_hd__xor2_1
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1097 final_adder.U$$182/B final_adder.U$$953/X VGND VGND VPWR VPWR
+ output355/A sky130_fd_sc_hd__xor2_1
XFILLER_113_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_50_3 dadda_fa_2_50_3/A dadda_fa_2_50_3/B dadda_fa_2_50_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/B dadda_fa_3_50_3/B sky130_fd_sc_hd__fa_1
XFILLER_22_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_43_2 U$$2753/X U$$2886/X input194/X VGND VGND VPWR VPWR dadda_fa_3_44_1/A
+ dadda_fa_3_43_3/A sky130_fd_sc_hd__fa_1
XFILLER_54_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3140 U$$3551/A1 U$$3148/A2 input121/X U$$3148/B2 VGND VGND VPWR VPWR U$$3141/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_20_1 dadda_fa_5_20_1/A dadda_fa_5_20_1/B dadda_fa_5_20_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_21_0/B dadda_fa_7_20_0/A sky130_fd_sc_hd__fa_1
XFILLER_19_471 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3151 U$$3151/A VGND VGND VPWR VPWR U$$3151/Y sky130_fd_sc_hd__inv_1
XU$$3162 U$$3162/A U$$3188/B VGND VGND VPWR VPWR U$$3162/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_36_1 U$$1143/X U$$1276/X U$$1409/X VGND VGND VPWR VPWR dadda_fa_3_37_0/CIN
+ dadda_fa_3_36_2/CIN sky130_fd_sc_hd__fa_1
XU$$3173 U$$842/B1 U$$3263/A2 input127/X U$$3263/B2 VGND VGND VPWR VPWR U$$3174/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_13_0 dadda_fa_5_13_0/A dadda_fa_5_13_0/B dadda_fa_5_13_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_14_0/A dadda_fa_6_13_0/CIN sky130_fd_sc_hd__fa_1
XU$$3184 U$$3184/A U$$3188/B VGND VGND VPWR VPWR U$$3184/X sky130_fd_sc_hd__xor2_1
XU$$3195 U$$727/B1 U$$3207/A2 U$$3606/B1 U$$3207/B2 VGND VGND VPWR VPWR U$$3196/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2450 U$$2450/A U$$2454/B VGND VGND VPWR VPWR U$$2450/X sky130_fd_sc_hd__xor2_1
XU$$2461 U$$3281/B1 U$$2463/A2 U$$3148/A1 U$$2463/B2 VGND VGND VPWR VPWR U$$2462/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_29_0 U$$65/X U$$198/X U$$331/X VGND VGND VPWR VPWR dadda_fa_3_30_1/B dadda_fa_3_29_3/A
+ sky130_fd_sc_hd__fa_1
XU$$2472 U$$2472/A1 U$$2524/A2 U$$2609/B1 U$$2524/B2 VGND VGND VPWR VPWR U$$2473/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2483 U$$2483/A U$$2491/B VGND VGND VPWR VPWR U$$2483/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2494 U$$3453/A1 U$$2524/A2 U$$3727/B1 U$$2524/B2 VGND VGND VPWR VPWR U$$2495/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1760 U$$2582/A1 U$$1764/A2 U$$527/B1 U$$1764/B2 VGND VGND VPWR VPWR U$$1761/A
+ sky130_fd_sc_hd__a22o_1
XU$$1771 U$$1771/A input18/X VGND VGND VPWR VPWR U$$1771/X sky130_fd_sc_hd__xor2_1
XFILLER_148_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1782 input19/X VGND VGND VPWR VPWR U$$1784/B sky130_fd_sc_hd__inv_1
XFILLER_194_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1793 U$$2065/B1 U$$1819/A2 U$$2343/A1 U$$1819/B2 VGND VGND VPWR VPWR U$$1794/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput70 b[14] VGND VGND VPWR VPWR input70/X sky130_fd_sc_hd__buf_6
Xinput81 b[24] VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_6
Xinput92 b[34] VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__buf_8
XFILLER_66_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_58_2 dadda_fa_4_58_2/A dadda_fa_4_58_2/B dadda_fa_4_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_59_0/CIN dadda_fa_5_58_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$401 final_adder.U$$400/B final_adder.U$$279/X final_adder.U$$275/X
+ VGND VGND VPWR VPWR final_adder.U$$401/X sky130_fd_sc_hd__a21o_1
XTAP_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$412 final_adder.U$$416/B final_adder.U$$412/B VGND VGND VPWR VPWR
+ final_adder.U$$536/B sky130_fd_sc_hd__and2_1
XTAP_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$423 final_adder.U$$422/B final_adder.U$$301/X final_adder.U$$297/X
+ VGND VGND VPWR VPWR final_adder.U$$423/X sky130_fd_sc_hd__a21o_1
XTAP_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$434 final_adder.U$$438/B final_adder.U$$434/B VGND VGND VPWR VPWR
+ final_adder.U$$558/B sky130_fd_sc_hd__and2_1
XFILLER_184_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$445 final_adder.U$$444/B final_adder.U$$323/X final_adder.U$$319/X
+ VGND VGND VPWR VPWR final_adder.U$$445/X sky130_fd_sc_hd__a21o_1
XTAP_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$456 final_adder.U$$460/B final_adder.U$$456/B VGND VGND VPWR VPWR
+ final_adder.U$$580/B sky130_fd_sc_hd__and2_1
XTAP_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater660 U$$805/B2 VGND VGND VPWR VPWR U$$759/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_7_28_0 dadda_fa_7_28_0/A dadda_fa_7_28_0/B dadda_fa_7_28_0/CIN VGND VGND
+ VPWR VPWR _325_/D _196_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$467 final_adder.U$$466/B final_adder.U$$345/X final_adder.U$$341/X
+ VGND VGND VPWR VPWR final_adder.U$$467/X sky130_fd_sc_hd__a21o_1
XU$$306 U$$717/A1 U$$316/A2 U$$34/A1 U$$316/B2 VGND VGND VPWR VPWR U$$307/A sky130_fd_sc_hd__a22o_1
XTAP_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater671 U$$4252/X VGND VGND VPWR VPWR U$$4297/B2 sky130_fd_sc_hd__buf_4
XFILLER_123_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$478 final_adder.U$$482/B final_adder.U$$478/B VGND VGND VPWR VPWR
+ final_adder.U$$602/B sky130_fd_sc_hd__and2_1
XTAP_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$317 U$$317/A U$$317/B VGND VGND VPWR VPWR U$$317/X sky130_fd_sc_hd__xor2_1
XFILLER_85_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater682 U$$521/B2 VGND VGND VPWR VPWR U$$515/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$489 final_adder.U$$488/B final_adder.U$$367/X final_adder.U$$363/X
+ VGND VGND VPWR VPWR final_adder.U$$489/X sky130_fd_sc_hd__a21o_1
XU$$328 U$$328/A1 U$$350/A2 U$$328/B1 U$$350/B2 VGND VGND VPWR VPWR U$$329/A sky130_fd_sc_hd__a22o_1
Xrepeater693 U$$4115/X VGND VGND VPWR VPWR U$$4240/B2 sky130_fd_sc_hd__buf_4
XFILLER_123_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$339 U$$339/A U$$343/B VGND VGND VPWR VPWR U$$339/X sky130_fd_sc_hd__xor2_1
XFILLER_198_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_636 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_674 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1206 U$$651/B VGND VGND VPWR VPWR U$$579/B sky130_fd_sc_hd__clkbuf_8
XFILLER_165_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1217 U$$504/B VGND VGND VPWR VPWR U$$474/B sky130_fd_sc_hd__buf_6
Xrepeater1228 U$$4366/B VGND VGND VPWR VPWR U$$4354/B sky130_fd_sc_hd__buf_4
XFILLER_148_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1239 input58/X VGND VGND VPWR VPWR U$$4247/A sky130_fd_sc_hd__buf_6
XFILLER_10_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_60_2 dadda_fa_3_60_2/A dadda_fa_3_60_2/B dadda_fa_3_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_1/A dadda_fa_4_60_2/B sky130_fd_sc_hd__fa_1
XFILLER_171_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_53_1 dadda_fa_3_53_1/A dadda_fa_3_53_1/B dadda_fa_3_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_0/CIN dadda_fa_4_53_2/A sky130_fd_sc_hd__fa_1
XFILLER_103_991 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_69_1 U$$810/X U$$943/X U$$1076/X VGND VGND VPWR VPWR dadda_fa_1_70_6/B
+ dadda_fa_1_69_8/A sky130_fd_sc_hd__fa_1
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_30_0 dadda_fa_6_30_0/A dadda_fa_6_30_0/B dadda_fa_6_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_31_0/B dadda_fa_7_30_0/CIN sky130_fd_sc_hd__fa_2
XTAP_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_46_0 dadda_fa_3_46_0/A dadda_fa_3_46_0/B dadda_fa_3_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_0/B dadda_fa_4_46_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_57_83 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$840 U$$18/A1 U$$872/A2 U$$979/A1 U$$872/B2 VGND VGND VPWR VPWR U$$841/A sky130_fd_sc_hd__a22o_1
XFILLER_1_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$851 U$$851/A U$$877/B VGND VGND VPWR VPWR U$$851/X sky130_fd_sc_hd__xor2_1
XFILLER_16_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$862 U$$997/B1 U$$882/A2 U$$864/A1 U$$882/B2 VGND VGND VPWR VPWR U$$863/A sky130_fd_sc_hd__a22o_1
XFILLER_91_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1001 U$$42/A1 U$$999/A2 U$$866/A1 U$$999/B2 VGND VGND VPWR VPWR U$$1002/A sky130_fd_sc_hd__a22o_1
XFILLER_32_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1012 U$$1012/A U$$998/B VGND VGND VPWR VPWR U$$1012/X sky130_fd_sc_hd__xor2_1
XFILLER_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$873 U$$873/A U$$877/B VGND VGND VPWR VPWR U$$873/X sky130_fd_sc_hd__xor2_1
XU$$884 U$$62/A1 U$$892/A2 U$$62/B1 U$$892/B2 VGND VGND VPWR VPWR U$$885/A sky130_fd_sc_hd__a22o_1
XU$$1023 U$$62/B1 U$$993/A2 U$$888/A1 U$$993/B2 VGND VGND VPWR VPWR U$$1024/A sky130_fd_sc_hd__a22o_1
XFILLER_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$895 U$$895/A U$$945/B VGND VGND VPWR VPWR U$$895/X sky130_fd_sc_hd__xor2_1
XFILLER_73_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1034 U$$1034/A U$$998/B VGND VGND VPWR VPWR U$$1034/X sky130_fd_sc_hd__xor2_1
XU$$1045 U$$84/B1 U$$965/A2 U$$910/A1 U$$965/B2 VGND VGND VPWR VPWR U$$1046/A sky130_fd_sc_hd__a22o_1
XFILLER_71_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1056 U$$1056/A U$$1084/B VGND VGND VPWR VPWR U$$1056/X sky130_fd_sc_hd__xor2_1
XU$$1067 U$$2709/B1 U$$963/X U$$2711/B1 U$$964/X VGND VGND VPWR VPWR U$$1068/A sky130_fd_sc_hd__a22o_1
XFILLER_32_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1078 U$$1078/A U$$1084/B VGND VGND VPWR VPWR U$$1078/X sky130_fd_sc_hd__xor2_1
XU$$1089 U$$952/A1 U$$1093/A2 U$$954/A1 U$$1093/B2 VGND VGND VPWR VPWR U$$1090/A sky130_fd_sc_hd__a22o_1
XFILLER_176_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_972 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_103_0 dadda_fa_7_103_0/A dadda_fa_7_103_0/B dadda_fa_7_103_0/CIN VGND
+ VGND VPWR VPWR _400_/D _271_/D sky130_fd_sc_hd__fa_1
XFILLER_8_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_98_3 U$$3528/X U$$3661/X U$$3794/X VGND VGND VPWR VPWR dadda_fa_3_99_1/CIN
+ dadda_fa_3_98_3/B sky130_fd_sc_hd__fa_1
XFILLER_176_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_68_1 dadda_fa_5_68_1/A dadda_fa_5_68_1/B dadda_fa_5_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_69_0/B dadda_fa_7_68_0/A sky130_fd_sc_hd__fa_1
XFILLER_98_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_107_0 U$$3013/Y U$$3147/X U$$3280/X VGND VGND VPWR VPWR dadda_fa_3_108_3/CIN
+ dadda_fa_4_107_0/A sky130_fd_sc_hd__fa_1
XFILLER_207_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_271 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2280 U$$2691/A1 U$$2316/A2 U$$3102/B1 U$$2316/B2 VGND VGND VPWR VPWR U$$2281/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2291 U$$2291/A U$$2317/B VGND VGND VPWR VPWR U$$2291/X sky130_fd_sc_hd__xor2_1
XFILLER_210_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1590 U$$1590/A U$$1592/B VGND VGND VPWR VPWR U$$1590/X sky130_fd_sc_hd__xor2_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1014 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_70_1 dadda_fa_4_70_1/A dadda_fa_4_70_1/B dadda_fa_4_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/B dadda_fa_5_70_1/B sky130_fd_sc_hd__fa_1
XFILLER_118_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_86_1 U$$1908/X U$$2041/X U$$2174/X VGND VGND VPWR VPWR dadda_fa_2_87_3/A
+ dadda_fa_2_86_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_63_0 dadda_fa_4_63_0/A dadda_fa_4_63_0/B dadda_fa_4_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/A dadda_fa_5_63_1/A sky130_fd_sc_hd__fa_1
XFILLER_89_466 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_79_0 U$$1095/Y U$$1229/X U$$1362/X VGND VGND VPWR VPWR dadda_fa_2_80_0/B
+ dadda_fa_2_79_3/B sky130_fd_sc_hd__fa_1
XFILLER_104_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$220 final_adder.U$$220/A final_adder.U$$220/B VGND VGND VPWR VPWR
+ final_adder.U$$348/B sky130_fd_sc_hd__and2_1
XTAP_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$231 final_adder.U$$230/B final_adder.U$$231/A2 final_adder.U$$231/B1
+ VGND VGND VPWR VPWR final_adder.U$$231/X sky130_fd_sc_hd__a21o_1
XTAP_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$242 final_adder.U$$242/A final_adder.U$$242/B VGND VGND VPWR VPWR
+ final_adder.U$$370/B sky130_fd_sc_hd__and2_1
XTAP_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3909 U$$3909/A U$$3909/B VGND VGND VPWR VPWR U$$3909/X sky130_fd_sc_hd__xor2_1
XTAP_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$253 final_adder.U$$3/SUM final_adder.U$$253/A2 final_adder.U$$3/COUT
+ VGND VGND VPWR VPWR final_adder.U$$253/X sky130_fd_sc_hd__a21o_1
XTAP_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$264 final_adder.U$$266/B final_adder.U$$264/B VGND VGND VPWR VPWR
+ final_adder.U$$390/B sky130_fd_sc_hd__and2_1
XTAP_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$103 U$$103/A U$$111/B VGND VGND VPWR VPWR U$$103/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$275 final_adder.U$$274/B final_adder.U$$149/X final_adder.U$$147/X
+ VGND VGND VPWR VPWR final_adder.U$$275/X sky130_fd_sc_hd__a21o_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$114 U$$251/A1 U$$122/A2 U$$116/A1 U$$122/B2 VGND VGND VPWR VPWR U$$115/A sky130_fd_sc_hd__a22o_1
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$286 final_adder.U$$288/B final_adder.U$$286/B VGND VGND VPWR VPWR
+ final_adder.U$$412/B sky130_fd_sc_hd__and2_1
Xrepeater490 U$$3388/A2 VGND VGND VPWR VPWR U$$3394/A2 sky130_fd_sc_hd__buf_4
XTAP_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$125 U$$125/A U$$127/B VGND VGND VPWR VPWR U$$125/X sky130_fd_sc_hd__xor2_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$297 final_adder.U$$296/B final_adder.U$$171/X final_adder.U$$169/X
+ VGND VGND VPWR VPWR final_adder.U$$297/X sky130_fd_sc_hd__a21o_1
XTAP_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$136 U$$136/A VGND VGND VPWR VPWR U$$136/Y sky130_fd_sc_hd__inv_1
XFILLER_45_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$147 U$$8/B1 U$$165/A2 U$$12/A1 U$$165/B2 VGND VGND VPWR VPWR U$$148/A sky130_fd_sc_hd__a22o_1
XFILLER_166_1228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$158 U$$158/A U$$160/B VGND VGND VPWR VPWR U$$158/X sky130_fd_sc_hd__xor2_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$169 U$$717/A1 U$$175/A2 U$$34/A1 U$$175/B2 VGND VGND VPWR VPWR U$$170/A sky130_fd_sc_hd__a22o_1
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_783 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1050 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_393_ _394_/CLK _393_/D VGND VGND VPWR VPWR _393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_1072 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1003 U$$3356/A1 VGND VGND VPWR VPWR U$$890/A1 sky130_fd_sc_hd__buf_4
XFILLER_86_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1014 input87/X VGND VGND VPWR VPWR U$$3300/A1 sky130_fd_sc_hd__buf_6
XFILLER_142_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1025 U$$3215/A1 VGND VGND VPWR VPWR U$$610/B1 sky130_fd_sc_hd__buf_4
Xrepeater1036 U$$3211/B1 VGND VGND VPWR VPWR U$$610/A1 sky130_fd_sc_hd__buf_8
Xdadda_fa_6_78_0 dadda_fa_6_78_0/A dadda_fa_6_78_0/B dadda_fa_6_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_79_0/B dadda_fa_7_78_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1047 input83/X VGND VGND VPWR VPWR U$$4442/B1 sky130_fd_sc_hd__buf_6
XFILLER_182_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1058 U$$330/A1 VGND VGND VPWR VPWR U$$328/B1 sky130_fd_sc_hd__buf_4
Xrepeater1069 U$$4027/A1 VGND VGND VPWR VPWR U$$874/B1 sky130_fd_sc_hd__buf_6
XFILLER_49_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$670 U$$807/A1 U$$552/X U$$807/B1 U$$553/X VGND VGND VPWR VPWR U$$671/A sky130_fd_sc_hd__a22o_1
XU$$681 U$$681/A U$$683/B VGND VGND VPWR VPWR U$$681/X sky130_fd_sc_hd__xor2_1
XFILLER_211_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$692 U$$692/A U$$712/B VGND VGND VPWR VPWR U$$692/X sky130_fd_sc_hd__xor2_1
XFILLER_204_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_394 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_80_0 dadda_fa_5_80_0/A dadda_fa_5_80_0/B dadda_fa_5_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_81_0/A dadda_fa_6_80_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_96_0 U$$2460/X U$$2593/X U$$2726/X VGND VGND VPWR VPWR dadda_fa_3_97_0/B
+ dadda_fa_3_96_2/B sky130_fd_sc_hd__fa_1
XFILLER_133_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1570 input116/X VGND VGND VPWR VPWR U$$4504/A1 sky130_fd_sc_hd__buf_4
Xrepeater1581 U$$2582/A1 VGND VGND VPWR VPWR U$$938/A1 sky130_fd_sc_hd__clkbuf_8
Xrepeater1592 U$$3813/A1 VGND VGND VPWR VPWR U$$251/A1 sky130_fd_sc_hd__buf_6
XFILLER_160_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_72_7 dadda_fa_1_72_7/A dadda_fa_1_72_7/B dadda_fa_1_72_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_73_2/CIN dadda_fa_2_72_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_65_6 dadda_fa_1_65_6/A dadda_fa_1_65_6/B dadda_fa_1_65_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_2/B dadda_fa_2_65_5/B sky130_fd_sc_hd__fa_1
XFILLER_104_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_5 U$$3581/X U$$3714/X U$$3847/X VGND VGND VPWR VPWR dadda_fa_2_59_2/A
+ dadda_fa_2_58_5/A sky130_fd_sc_hd__fa_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_95_0 dadda_fa_7_95_0/A dadda_fa_7_95_0/B dadda_fa_7_95_0/CIN VGND VGND
+ VPWR VPWR _392_/D _263_/D sky130_fd_sc_hd__fa_2
XFILLER_202_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_780 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_666 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$417_1762 VGND VGND VPWR VPWR U$$417_1762/HI U$$417/A1 sky130_fd_sc_hd__conb_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4407 U$$4407/A U$$4407/B VGND VGND VPWR VPWR U$$4407/X sky130_fd_sc_hd__xor2_1
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4418 U$$4418/A1 U$$4388/X U$$4420/A1 U$$4426/B2 VGND VGND VPWR VPWR U$$4419/A
+ sky130_fd_sc_hd__a22o_1
XU$$4429 U$$4429/A U$$4429/B VGND VGND VPWR VPWR U$$4429/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_110_0 dadda_fa_6_110_0/A dadda_fa_6_110_0/B dadda_fa_6_110_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_111_0/B dadda_fa_7_110_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3706 U$$3706/A U$$3794/B VGND VGND VPWR VPWR U$$3706/X sky130_fd_sc_hd__xor2_1
XTAP_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3717 U$$3852/B1 U$$3753/A2 U$$3719/A1 U$$3753/B2 VGND VGND VPWR VPWR U$$3718/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3728 U$$3728/A U$$3740/B VGND VGND VPWR VPWR U$$3728/X sky130_fd_sc_hd__xor2_1
XU$$3739 U$$4424/A1 U$$3739/A2 U$$3876/B1 U$$3739/B2 VGND VGND VPWR VPWR U$$3740/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_30_3 dadda_fa_3_30_3/A dadda_fa_3_30_3/B dadda_fa_3_30_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_31_1/B dadda_fa_4_30_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_23_2 U$$1117/X U$$1250/X U$$1383/X VGND VGND VPWR VPWR dadda_fa_4_24_1/A
+ dadda_fa_4_23_2/B sky130_fd_sc_hd__fa_1
XTAP_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_861 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_376_ _376_/CLK _376_/D VGND VGND VPWR VPWR _376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_75_5 dadda_fa_2_75_5/A dadda_fa_2_75_5/B dadda_fa_2_75_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_76_2/A dadda_fa_4_75_0/A sky130_fd_sc_hd__fa_1
XFILLER_123_861 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_68_4 dadda_fa_2_68_4/A dadda_fa_2_68_4/B dadda_fa_2_68_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_1/CIN dadda_fa_3_68_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_205_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_992 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1102_1711 VGND VGND VPWR VPWR U$$1102_1711/HI U$$1102/A1 sky130_fd_sc_hd__conb_1
XFILLER_192_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_105_1 dadda_fa_5_105_1/A dadda_fa_5_105_1/B dadda_fa_5_105_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_106_0/B dadda_fa_7_105_0/A sky130_fd_sc_hd__fa_1
XFILLER_121_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_70_4 U$$3871/X U$$4004/X U$$4137/X VGND VGND VPWR VPWR dadda_fa_2_71_1/CIN
+ dadda_fa_2_70_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_63_3 U$$3591/X U$$3724/X U$$3857/X VGND VGND VPWR VPWR dadda_fa_2_64_1/B
+ dadda_fa_2_63_4/B sky130_fd_sc_hd__fa_1
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_40_2 dadda_fa_4_40_2/A dadda_fa_4_40_2/B dadda_fa_4_40_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_41_0/CIN dadda_fa_5_40_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_56_2 U$$1981/X U$$2114/X U$$2247/X VGND VGND VPWR VPWR dadda_fa_2_57_1/A
+ dadda_fa_2_56_4/A sky130_fd_sc_hd__fa_1
XFILLER_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_33_1 dadda_fa_4_33_1/A dadda_fa_4_33_1/B dadda_fa_4_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/B dadda_fa_5_33_1/B sky130_fd_sc_hd__fa_1
XFILLER_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_49_1 U$$504/X U$$637/X U$$770/X VGND VGND VPWR VPWR dadda_fa_2_50_1/A
+ dadda_fa_2_49_4/A sky130_fd_sc_hd__fa_1
XFILLER_131_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_10_0 dadda_fa_7_10_0/A dadda_fa_7_10_0/B dadda_fa_7_10_0/CIN VGND VGND
+ VPWR VPWR _307_/D _178_/D sky130_fd_sc_hd__fa_1
XFILLER_131_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_26_0 dadda_fa_4_26_0/A dadda_fa_4_26_0/B dadda_fa_4_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/A dadda_fa_5_26_1/A sky130_fd_sc_hd__fa_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_230_ _359_/CLK _230_/D VGND VGND VPWR VPWR _230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_842 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_78_3 dadda_fa_3_78_3/A dadda_fa_3_78_3/B dadda_fa_3_78_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_79_1/B dadda_fa_4_78_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1076 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4204 input102/X U$$4226/A2 input103/X U$$4226/B2 VGND VGND VPWR VPWR U$$4205/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4215 U$$4215/A U$$4227/B VGND VGND VPWR VPWR U$$4215/X sky130_fd_sc_hd__xor2_1
XFILLER_120_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4226 U$$4361/B1 U$$4226/A2 U$$4228/A1 U$$4226/B2 VGND VGND VPWR VPWR U$$4227/A
+ sky130_fd_sc_hd__a22o_1
XU$$4237 U$$4237/A U$$4239/B VGND VGND VPWR VPWR U$$4237/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_15_0 U$$37/X U$$170/X VGND VGND VPWR VPWR dadda_fa_4_16_2/A dadda_ha_3_15_0/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_20_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3503 U$$3775/B1 U$$3503/A2 U$$3642/A1 U$$3503/B2 VGND VGND VPWR VPWR U$$3504/A
+ sky130_fd_sc_hd__a22o_1
XU$$4248 input59/X VGND VGND VPWR VPWR U$$4250/B sky130_fd_sc_hd__inv_1
XFILLER_168_1109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3514 U$$3514/A U$$3518/B VGND VGND VPWR VPWR U$$3514/X sky130_fd_sc_hd__xor2_1
XU$$4259 U$$4396/A1 U$$4275/A2 U$$4398/A1 U$$4275/B2 VGND VGND VPWR VPWR U$$4260/A
+ sky130_fd_sc_hd__a22o_1
XU$$1641_1720 VGND VGND VPWR VPWR U$$1641_1720/HI U$$1641/B1 sky130_fd_sc_hd__conb_1
XU$$3525 U$$4210/A1 U$$3527/A2 U$$4210/B1 U$$3527/B2 VGND VGND VPWR VPWR U$$3526/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3536 U$$3536/A U$$3561/A VGND VGND VPWR VPWR U$$3536/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2802 U$$3211/B1 U$$2810/A2 U$$3352/A1 U$$2810/B2 VGND VGND VPWR VPWR U$$2803/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3547 U$$122/A1 U$$3549/A2 U$$3547/B1 U$$3549/B2 VGND VGND VPWR VPWR U$$3548/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3558 U$$3558/A U$$3561/A VGND VGND VPWR VPWR U$$3558/X sky130_fd_sc_hd__xor2_1
XFILLER_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2813 U$$2813/A U$$2825/B VGND VGND VPWR VPWR U$$2813/X sky130_fd_sc_hd__xor2_1
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3569 U$$3569/A U$$3609/B VGND VGND VPWR VPWR U$$3569/X sky130_fd_sc_hd__xor2_1
XFILLER_45_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2824 U$$3646/A1 U$$2828/A2 U$$4468/B1 U$$2828/B2 VGND VGND VPWR VPWR U$$2825/A
+ sky130_fd_sc_hd__a22o_1
XU$$2835 U$$2835/A U$$2837/B VGND VGND VPWR VPWR U$$2835/X sky130_fd_sc_hd__xor2_1
XFILLER_61_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2846 U$$2981/B1 U$$2874/A2 U$$4492/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2847/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2857 U$$2857/A U$$2869/B VGND VGND VPWR VPWR U$$2857/X sky130_fd_sc_hd__xor2_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 U$$3082/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_206_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2868 U$$3414/B1 U$$2868/A2 U$$3281/A1 U$$2868/B2 VGND VGND VPWR VPWR U$$2869/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 U$$3227/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_162 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2879 input38/X VGND VGND VPWR VPWR U$$2879/Y sky130_fd_sc_hd__inv_1
XANTENNA_173 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_184 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1014 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4407_1780 VGND VGND VPWR VPWR U$$4407_1780/HI U$$4407/B sky130_fd_sc_hd__conb_1
XFILLER_42_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_359_ _359_/CLK _359_/D VGND VGND VPWR VPWR _359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_750 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_80_3 dadda_fa_2_80_3/A dadda_fa_2_80_3/B dadda_fa_2_80_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/B dadda_fa_3_80_3/B sky130_fd_sc_hd__fa_1
XFILLER_103_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_73_2 dadda_fa_2_73_2/A dadda_fa_2_73_2/B dadda_fa_2_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/A dadda_fa_3_73_3/A sky130_fd_sc_hd__fa_1
XFILLER_155_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_222 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_50_1 dadda_fa_5_50_1/A dadda_fa_5_50_1/B dadda_fa_5_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_51_0/B dadda_fa_7_50_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_66_1 dadda_fa_2_66_1/A dadda_fa_2_66_1/B dadda_fa_2_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_0/CIN dadda_fa_3_66_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$819 final_adder.U$$786/A final_adder.U$$619/X final_adder.U$$707/X
+ VGND VGND VPWR VPWR final_adder.U$$819/X sky130_fd_sc_hd__a21o_1
XFILLER_151_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_43_0 dadda_fa_5_43_0/A dadda_fa_5_43_0/B dadda_fa_5_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_44_0/A dadda_fa_6_43_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_59_0 dadda_fa_2_59_0/A dadda_fa_2_59_0/B dadda_fa_2_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_0/B dadda_fa_3_59_2/B sky130_fd_sc_hd__fa_1
XFILLER_111_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 a[10] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_2
XFILLER_84_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$0 _296_/Q _168_/Q VGND VGND VPWR VPWR final_adder.U$$255/A2 final_adder.U$$0/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_69_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_934 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_88_2 dadda_fa_4_88_2/A dadda_fa_4_88_2/B dadda_fa_4_88_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_89_0/CIN dadda_fa_5_88_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_156_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput350 output350/A VGND VGND VPWR VPWR o[69] sky130_fd_sc_hd__buf_2
Xoutput361 output361/A VGND VGND VPWR VPWR o[79] sky130_fd_sc_hd__buf_2
Xdadda_fa_7_58_0 dadda_fa_7_58_0/A dadda_fa_7_58_0/B dadda_fa_7_58_0/CIN VGND VGND
+ VPWR VPWR _355_/D _226_/D sky130_fd_sc_hd__fa_1
XFILLER_121_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput372 output372/A VGND VGND VPWR VPWR o[89] sky130_fd_sc_hd__buf_2
XFILLER_0_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput383 output383/A VGND VGND VPWR VPWR o[99] sky130_fd_sc_hd__buf_2
XFILLER_82_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_61_0 U$$1991/X U$$2124/X U$$2257/X VGND VGND VPWR VPWR dadda_fa_2_62_0/B
+ dadda_fa_2_61_3/B sky130_fd_sc_hd__fa_1
XFILLER_75_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2109 U$$3614/B1 U$$2113/A2 U$$3481/A1 U$$2113/B2 VGND VGND VPWR VPWR U$$2110/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1408 U$$721/B1 U$$1434/A2 U$$997/B1 U$$1434/B2 VGND VGND VPWR VPWR U$$1409/A sky130_fd_sc_hd__a22o_1
XU$$1419 U$$1419/A U$$1423/B VGND VGND VPWR VPWR U$$1419/X sky130_fd_sc_hd__xor2_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1003 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_213_ _342_/CLK _213_/D VGND VGND VPWR VPWR _213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_90_2 dadda_fa_3_90_2/A dadda_fa_3_90_2/B dadda_fa_3_90_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_1/A dadda_fa_4_90_2/B sky130_fd_sc_hd__fa_2
XFILLER_164_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1097 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_83_1 dadda_fa_3_83_1/A dadda_fa_3_83_1/B dadda_fa_3_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_0/CIN dadda_fa_4_83_2/A sky130_fd_sc_hd__fa_1
XFILLER_152_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_60_0 dadda_fa_6_60_0/A dadda_fa_6_60_0/B dadda_fa_6_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_61_0/B dadda_fa_7_60_0/CIN sky130_fd_sc_hd__fa_1
XU$$4437_1795 VGND VGND VPWR VPWR U$$4437_1795/HI U$$4437/B sky130_fd_sc_hd__conb_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_76_0 dadda_fa_3_76_0/A dadda_fa_3_76_0/B dadda_fa_3_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_0/B dadda_fa_4_76_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4001 U$$4273/B1 U$$4035/A2 U$$4275/B1 U$$4035/B2 VGND VGND VPWR VPWR U$$4002/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4012 U$$4012/A U$$4012/B VGND VGND VPWR VPWR U$$4012/X sky130_fd_sc_hd__xor2_1
XU$$4023 input78/X U$$4043/A2 input79/X U$$4043/B2 VGND VGND VPWR VPWR U$$4024/A sky130_fd_sc_hd__a22o_1
XU$$4034 U$$4034/A U$$4036/B VGND VGND VPWR VPWR U$$4034/X sky130_fd_sc_hd__xor2_1
XFILLER_65_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4045 U$$4045/A1 U$$4107/A2 input91/X U$$4107/B2 VGND VGND VPWR VPWR U$$4046/A
+ sky130_fd_sc_hd__a22o_1
XU$$3300 U$$3300/A1 U$$3320/A2 U$$3300/B1 U$$3320/B2 VGND VGND VPWR VPWR U$$3301/A
+ sky130_fd_sc_hd__a22o_1
XU$$3311 U$$3311/A U$$3395/B VGND VGND VPWR VPWR U$$3311/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_1 dadda_fa_4_112_1/A dadda_fa_4_112_1/B dadda_fa_4_112_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_113_0/B dadda_fa_5_112_1/B sky130_fd_sc_hd__fa_1
XU$$4056 U$$4056/A U$$4080/B VGND VGND VPWR VPWR U$$4056/X sky130_fd_sc_hd__xor2_1
XFILLER_24_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4067 U$$4476/B1 U$$4077/A2 U$$4343/A1 U$$4077/B2 VGND VGND VPWR VPWR U$$4068/A
+ sky130_fd_sc_hd__a22o_1
XU$$3322 U$$4005/B1 U$$3348/A2 U$$4009/A1 U$$3346/B2 VGND VGND VPWR VPWR U$$3323/A
+ sky130_fd_sc_hd__a22o_1
XU$$4078 U$$4078/A U$$4078/B VGND VGND VPWR VPWR U$$4078/X sky130_fd_sc_hd__xor2_1
XU$$3333 U$$3333/A U$$3375/B VGND VGND VPWR VPWR U$$3333/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4089 U$$4361/B1 U$$4101/A2 U$$4228/A1 U$$4101/B2 VGND VGND VPWR VPWR U$$4090/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3344 U$$3344/A1 U$$3378/A2 U$$741/B1 U$$3346/B2 VGND VGND VPWR VPWR U$$3345/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2610 U$$2610/A U$$2624/B VGND VGND VPWR VPWR U$$2610/X sky130_fd_sc_hd__xor2_1
XFILLER_62_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3355 U$$3355/A U$$3389/B VGND VGND VPWR VPWR U$$3355/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_105_0 dadda_fa_4_105_0/A dadda_fa_4_105_0/B dadda_fa_4_105_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/A dadda_fa_5_105_1/A sky130_fd_sc_hd__fa_1
XFILLER_34_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2621 U$$2621/A1 U$$2625/A2 U$$2623/A1 U$$2625/B2 VGND VGND VPWR VPWR U$$2622/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_38_5 dadda_fa_2_38_5/A dadda_fa_2_38_5/B dadda_fa_2_38_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_39_2/A dadda_fa_4_38_0/A sky130_fd_sc_hd__fa_1
XFILLER_74_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3366 U$$3366/A1 U$$3292/X U$$3366/B1 U$$3293/X VGND VGND VPWR VPWR U$$3367/A sky130_fd_sc_hd__a22o_1
XFILLER_206_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3377 U$$3377/A U$$3377/B VGND VGND VPWR VPWR U$$3377/X sky130_fd_sc_hd__xor2_1
XU$$2632 U$$2632/A U$$2650/B VGND VGND VPWR VPWR U$$2632/X sky130_fd_sc_hd__xor2_1
XU$$2643 U$$38/B1 U$$2727/A2 U$$4013/B1 U$$2727/B2 VGND VGND VPWR VPWR U$$2644/A sky130_fd_sc_hd__a22o_1
XU$$3388 U$$783/B1 U$$3388/A2 U$$650/A1 U$$3390/B2 VGND VGND VPWR VPWR U$$3389/A sky130_fd_sc_hd__a22o_1
XU$$3399 U$$3399/A U$$3417/B VGND VGND VPWR VPWR U$$3399/X sky130_fd_sc_hd__xor2_1
XFILLER_179_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2654 U$$2654/A U$$2658/B VGND VGND VPWR VPWR U$$2654/X sky130_fd_sc_hd__xor2_1
XFILLER_94_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2665 U$$4309/A1 U$$2607/X U$$4309/B1 U$$2608/X VGND VGND VPWR VPWR U$$2666/A sky130_fd_sc_hd__a22o_1
XU$$1920 input22/X VGND VGND VPWR VPWR U$$1920/Y sky130_fd_sc_hd__inv_1
XFILLER_55_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1931 U$$1931/A U$$1991/B VGND VGND VPWR VPWR U$$1931/X sky130_fd_sc_hd__xor2_1
XU$$2676 U$$2676/A U$$2680/B VGND VGND VPWR VPWR U$$2676/X sky130_fd_sc_hd__xor2_1
XU$$1942 U$$3584/B1 U$$1990/A2 U$$2901/B1 U$$1990/B2 VGND VGND VPWR VPWR U$$1943/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2687 U$$3646/A1 U$$2735/A2 U$$3922/A1 U$$2735/B2 VGND VGND VPWR VPWR U$$2688/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1953 U$$1953/A U$$1993/B VGND VGND VPWR VPWR U$$1953/X sky130_fd_sc_hd__xor2_1
XFILLER_34_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2698 U$$2698/A U$$2716/B VGND VGND VPWR VPWR U$$2698/X sky130_fd_sc_hd__xor2_1
XU$$1964 U$$44/B1 U$$1990/A2 U$$3747/A1 U$$1990/B2 VGND VGND VPWR VPWR U$$1965/A sky130_fd_sc_hd__a22o_1
XU$$1975 U$$1975/A U$$2017/B VGND VGND VPWR VPWR U$$1975/X sky130_fd_sc_hd__xor2_1
XFILLER_194_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1986 U$$2123/A1 U$$2016/A2 U$$616/B1 U$$2016/B2 VGND VGND VPWR VPWR U$$1987/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1997 U$$1997/A U$$2043/B VGND VGND VPWR VPWR U$$1997/X sky130_fd_sc_hd__xor2_1
XFILLER_14_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_98_1 dadda_fa_5_98_1/A dadda_fa_5_98_1/B dadda_fa_5_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_99_0/B dadda_fa_7_98_0/A sky130_fd_sc_hd__fa_1
XFILLER_135_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$605 final_adder.U$$604/B final_adder.U$$489/X final_adder.U$$481/X
+ VGND VGND VPWR VPWR final_adder.U$$605/X sky130_fd_sc_hd__a21o_1
XFILLER_84_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$616 final_adder.U$$616/A final_adder.U$$616/B VGND VGND VPWR VPWR
+ final_adder.U$$720/A sky130_fd_sc_hd__and2_1
Xrepeater820 U$$2060/X VGND VGND VPWR VPWR U$$2183/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater831 U$$1831/B2 VGND VGND VPWR VPWR U$$1839/B2 sky130_fd_sc_hd__buf_6
XFILLER_99_1025 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$638 final_adder.U$$654/B final_adder.U$$638/B VGND VGND VPWR VPWR
+ final_adder.U$$750/B sky130_fd_sc_hd__and2_1
XTAP_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater842 U$$1750/B2 VGND VGND VPWR VPWR U$$1706/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$649 final_adder.U$$648/B final_adder.U$$545/X final_adder.U$$529/X
+ VGND VGND VPWR VPWR final_adder.U$$649/X sky130_fd_sc_hd__a21o_1
Xrepeater853 U$$1512/X VGND VGND VPWR VPWR U$$1607/B2 sky130_fd_sc_hd__buf_6
XFILLER_38_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater864 U$$1504/B2 VGND VGND VPWR VPWR U$$1502/B2 sky130_fd_sc_hd__buf_6
Xrepeater875 U$$1281/B2 VGND VGND VPWR VPWR U$$1271/B2 sky130_fd_sc_hd__clkbuf_4
Xrepeater886 U$$1101/X VGND VGND VPWR VPWR U$$1204/B2 sky130_fd_sc_hd__buf_8
XFILLER_84_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater897 U$$4389/X VGND VGND VPWR VPWR U$$4432/B2 sky130_fd_sc_hd__buf_4
XFILLER_84_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$60 U$$60/A1 U$$94/A2 U$$62/A1 U$$94/B2 VGND VGND VPWR VPWR U$$61/A sky130_fd_sc_hd__a22o_1
XU$$71 U$$71/A U$$81/B VGND VGND VPWR VPWR U$$71/X sky130_fd_sc_hd__xor2_1
XU$$82 U$$82/A1 U$$98/A2 U$$84/A1 U$$98/B2 VGND VGND VPWR VPWR U$$83/A sky130_fd_sc_hd__a22o_1
XU$$93 U$$93/A U$$99/B VGND VGND VPWR VPWR U$$93/X sky130_fd_sc_hd__xor2_1
XFILLER_53_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_40 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_51 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _342_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_73 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_84 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_93_0 dadda_fa_4_93_0/A dadda_fa_4_93_0/B dadda_fa_4_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/A dadda_fa_5_93_1/A sky130_fd_sc_hd__fa_1
XANTENNA_95 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_107_2 U$$4211/X U$$4344/X U$$4477/X VGND VGND VPWR VPWR dadda_fa_4_108_1/A
+ dadda_fa_4_107_2/B sky130_fd_sc_hd__fa_1
XFILLER_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_984 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1205 U$$1205/A U$$1205/B VGND VGND VPWR VPWR U$$1205/X sky130_fd_sc_hd__xor2_1
XU$$1216 U$$942/A1 U$$1222/A2 U$$944/A1 U$$1222/B2 VGND VGND VPWR VPWR U$$1217/A sky130_fd_sc_hd__a22o_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1227 U$$1227/A U$$1232/A VGND VGND VPWR VPWR U$$1227/X sky130_fd_sc_hd__xor2_1
XFILLER_203_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1238 U$$1236/B input9/X input10/X U$$1233/Y VGND VGND VPWR VPWR U$$1238/X sky130_fd_sc_hd__a22o_2
XFILLER_206_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1249 U$$2206/B1 U$$1271/A2 U$$3032/A1 U$$1271/B2 VGND VGND VPWR VPWR U$$1250/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1376_1716 VGND VGND VPWR VPWR U$$1376_1716/HI U$$1376/A1 sky130_fd_sc_hd__conb_1
XFILLER_168_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1021 final_adder.U$$4/SUM final_adder.U$$381/X final_adder.U$$4/COUT
+ VGND VGND VPWR VPWR final_adder.U$$1029/B sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$1032 final_adder.U$$8/SUM final_adder.U$$503/X VGND VGND VPWR VPWR
+ output373/A sky130_fd_sc_hd__xor2_1
XFILLER_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1043 final_adder.U$$236/B final_adder.U$$1043/B VGND VGND VPWR VPWR
+ output295/A sky130_fd_sc_hd__xor2_1
XFILLER_156_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1054 final_adder.U$$224/A final_adder.U$$725/X VGND VGND VPWR VPWR
+ output308/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1065 final_adder.U$$214/B final_adder.U$$985/X VGND VGND VPWR VPWR
+ output320/A sky130_fd_sc_hd__xor2_1
XFILLER_171_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1076 final_adder.U$$202/A final_adder.U$$815/X VGND VGND VPWR VPWR
+ output332/A sky130_fd_sc_hd__xor2_1
XFILLER_194_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1087 final_adder.U$$192/B final_adder.U$$963/X VGND VGND VPWR VPWR
+ output344/A sky130_fd_sc_hd__xor2_1
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1098 final_adder.U$$180/A final_adder.U$$889/X VGND VGND VPWR VPWR
+ output356/A sky130_fd_sc_hd__xor2_1
XFILLER_194_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_50_4 dadda_fa_2_50_4/A dadda_fa_2_50_4/B dadda_fa_2_50_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_1/CIN dadda_fa_3_50_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2335_1731 VGND VGND VPWR VPWR U$$2335_1731/HI U$$2335/A1 sky130_fd_sc_hd__conb_1
Xdadda_fa_2_43_3 dadda_fa_2_43_3/A dadda_fa_2_43_3/B dadda_fa_2_43_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_1/B dadda_fa_3_43_3/B sky130_fd_sc_hd__fa_1
XU$$3130 U$$116/A1 U$$3132/A2 U$$3680/A1 U$$3132/B2 VGND VGND VPWR VPWR U$$3131/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3141 U$$3141/A U$$3150/A VGND VGND VPWR VPWR U$$3141/X sky130_fd_sc_hd__xor2_1
XFILLER_35_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3152 input41/X VGND VGND VPWR VPWR U$$3154/B sky130_fd_sc_hd__inv_1
XFILLER_19_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_36_2 U$$1542/X U$$1675/X U$$1808/X VGND VGND VPWR VPWR dadda_fa_3_37_1/A
+ dadda_fa_3_36_3/A sky130_fd_sc_hd__fa_1
XU$$3163 U$$3300/A1 U$$3187/A2 U$$3300/B1 U$$3187/B2 VGND VGND VPWR VPWR U$$3164/A
+ sky130_fd_sc_hd__a22o_1
XU$$3174 U$$3174/A U$$3264/B VGND VGND VPWR VPWR U$$3174/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2440 U$$2440/A U$$2466/A VGND VGND VPWR VPWR U$$2440/X sky130_fd_sc_hd__xor2_1
XFILLER_62_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3185 U$$4144/A1 U$$3187/A2 U$$4144/B1 U$$3187/B2 VGND VGND VPWR VPWR U$$3186/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_13_1 dadda_fa_5_13_1/A dadda_fa_5_13_1/B dadda_ha_4_13_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_14_0/B dadda_fa_7_13_0/A sky130_fd_sc_hd__fa_1
XFILLER_207_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2451 U$$4095/A1 U$$2459/A2 U$$3960/A1 U$$2459/B2 VGND VGND VPWR VPWR U$$2452/A
+ sky130_fd_sc_hd__a22o_1
XU$$3196 U$$3196/A U$$3208/B VGND VGND VPWR VPWR U$$3196/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_29_1 U$$464/X U$$597/X U$$730/X VGND VGND VPWR VPWR dadda_fa_3_30_1/CIN
+ dadda_fa_3_29_3/B sky130_fd_sc_hd__fa_1
XU$$2462 U$$2462/A U$$2465/A VGND VGND VPWR VPWR U$$2462/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2473 U$$2473/A U$$2525/B VGND VGND VPWR VPWR U$$2473/X sky130_fd_sc_hd__xor2_1
XU$$2484 U$$2621/A1 U$$2490/A2 U$$2623/A1 U$$2490/B2 VGND VGND VPWR VPWR U$$2485/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2495 U$$2495/A U$$2525/B VGND VGND VPWR VPWR U$$2495/X sky130_fd_sc_hd__xor2_1
XU$$1750 U$$928/A1 U$$1750/A2 U$$930/A1 U$$1750/B2 VGND VGND VPWR VPWR U$$1751/A sky130_fd_sc_hd__a22o_1
XFILLER_34_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1761 U$$1761/A U$$1765/B VGND VGND VPWR VPWR U$$1761/X sky130_fd_sc_hd__xor2_1
XFILLER_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_727 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1772 U$$2044/B1 U$$1648/X U$$4514/A1 U$$1649/X VGND VGND VPWR VPWR U$$1773/A sky130_fd_sc_hd__a22o_1
XFILLER_72_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1783 U$$1912/B VGND VGND VPWR VPWR U$$1783/Y sky130_fd_sc_hd__inv_1
XU$$1794 U$$1794/A U$$1820/B VGND VGND VPWR VPWR U$$1794/X sky130_fd_sc_hd__xor2_1
XFILLER_148_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput60 a[63] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_6
Xinput71 b[15] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__buf_12
Xinput82 b[25] VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__buf_6
Xinput93 b[35] VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__buf_8
XFILLER_66_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$402 final_adder.U$$406/B final_adder.U$$402/B VGND VGND VPWR VPWR
+ final_adder.U$$526/B sky130_fd_sc_hd__and2_1
XTAP_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$413 final_adder.U$$412/B final_adder.U$$291/X final_adder.U$$287/X
+ VGND VGND VPWR VPWR final_adder.U$$413/X sky130_fd_sc_hd__a21o_1
XTAP_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$424 final_adder.U$$428/B final_adder.U$$424/B VGND VGND VPWR VPWR
+ final_adder.U$$548/B sky130_fd_sc_hd__and2_1
XFILLER_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$435 final_adder.U$$434/B final_adder.U$$313/X final_adder.U$$309/X
+ VGND VGND VPWR VPWR final_adder.U$$435/X sky130_fd_sc_hd__a21o_1
XTAP_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$0_1709 VGND VGND VPWR VPWR U$$0_1709/HI U$$0/A sky130_fd_sc_hd__conb_1
Xfinal_adder.U$$446 final_adder.U$$450/B final_adder.U$$446/B VGND VGND VPWR VPWR
+ final_adder.U$$570/B sky130_fd_sc_hd__and2_1
XTAP_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater650 U$$938/B2 VGND VGND VPWR VPWR U$$892/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$457 final_adder.U$$456/B final_adder.U$$335/X final_adder.U$$331/X
+ VGND VGND VPWR VPWR final_adder.U$$457/X sky130_fd_sc_hd__a21o_1
XTAP_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater661 U$$690/X VGND VGND VPWR VPWR U$$805/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$468 final_adder.U$$472/B final_adder.U$$468/B VGND VGND VPWR VPWR
+ final_adder.U$$592/B sky130_fd_sc_hd__and2_1
XU$$307 U$$307/A U$$317/B VGND VGND VPWR VPWR U$$307/X sky130_fd_sc_hd__xor2_1
XTAP_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater672 U$$4252/X VGND VGND VPWR VPWR U$$4381/B2 sky130_fd_sc_hd__clkbuf_8
Xfinal_adder.U$$479 final_adder.U$$478/B final_adder.U$$357/X final_adder.U$$353/X
+ VGND VGND VPWR VPWR final_adder.U$$479/X sky130_fd_sc_hd__a21o_1
Xrepeater683 U$$527/B2 VGND VGND VPWR VPWR U$$521/B2 sky130_fd_sc_hd__buf_6
XU$$318 U$$44/A1 U$$340/A2 U$$46/A1 U$$340/B2 VGND VGND VPWR VPWR U$$319/A sky130_fd_sc_hd__a22o_1
XU$$329 U$$329/A U$$351/B VGND VGND VPWR VPWR U$$329/X sky130_fd_sc_hd__xor2_1
Xrepeater694 U$$4043/B2 VGND VGND VPWR VPWR U$$4011/B2 sky130_fd_sc_hd__buf_4
XFILLER_84_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_112_0 dadda_fa_3_112_0/A U$$3423/X U$$3556/X VGND VGND VPWR VPWR dadda_fa_4_113_1/B
+ dadda_fa_4_112_2/A sky130_fd_sc_hd__fa_1
Xrepeater1207 U$$684/A VGND VGND VPWR VPWR U$$651/B sky130_fd_sc_hd__buf_6
XU$$2874_1740 VGND VGND VPWR VPWR U$$2874_1740/HI U$$2874/B1 sky130_fd_sc_hd__conb_1
Xrepeater1218 U$$516/B VGND VGND VPWR VPWR U$$436/B sky130_fd_sc_hd__buf_4
XFILLER_10_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1229 U$$4370/B VGND VGND VPWR VPWR U$$4366/B sky130_fd_sc_hd__buf_8
XFILLER_49_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1252 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_60_3 dadda_fa_3_60_3/A dadda_fa_3_60_3/B dadda_fa_3_60_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_61_1/B dadda_fa_4_60_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_53_2 dadda_fa_3_53_2/A dadda_fa_3_53_2/B dadda_fa_3_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_1/A dadda_fa_4_53_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_0_69_2 U$$1209/X U$$1342/X U$$1475/X VGND VGND VPWR VPWR dadda_fa_1_70_6/CIN
+ dadda_fa_1_69_8/B sky130_fd_sc_hd__fa_1
XFILLER_75_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_46_1 dadda_fa_3_46_1/A dadda_fa_3_46_1/B dadda_fa_3_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_0/CIN dadda_fa_4_46_2/A sky130_fd_sc_hd__fa_1
XTAP_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_23_0 dadda_fa_6_23_0/A dadda_fa_6_23_0/B dadda_fa_6_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_24_0/B dadda_fa_7_23_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_21_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_39_0 dadda_fa_3_39_0/A dadda_fa_3_39_0/B dadda_fa_3_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_0/B dadda_fa_4_39_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$991 final_adder.U$$220/A final_adder.U$$833/X final_adder.U$$991/B1
+ VGND VGND VPWR VPWR final_adder.U$$991/X sky130_fd_sc_hd__a21o_1
XU$$830 U$$967/A1 U$$918/A2 U$$832/A1 U$$918/B2 VGND VGND VPWR VPWR U$$831/A sky130_fd_sc_hd__a22o_1
XU$$841 U$$841/A U$$847/B VGND VGND VPWR VPWR U$$841/X sky130_fd_sc_hd__xor2_1
XFILLER_44_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$852 U$$987/B1 U$$872/A2 U$$854/A1 U$$872/B2 VGND VGND VPWR VPWR U$$853/A sky130_fd_sc_hd__a22o_1
XU$$863 U$$863/A U$$883/B VGND VGND VPWR VPWR U$$863/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1002 U$$1002/A U$$996/B VGND VGND VPWR VPWR U$$1002/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1013 U$$54/A1 U$$997/A2 U$$330/A1 U$$997/B2 VGND VGND VPWR VPWR U$$1014/A sky130_fd_sc_hd__a22o_1
XU$$874 U$$52/A1 U$$906/A2 U$$874/B1 U$$906/B2 VGND VGND VPWR VPWR U$$875/A sky130_fd_sc_hd__a22o_1
XU$$1024 U$$1024/A U$$994/B VGND VGND VPWR VPWR U$$1024/X sky130_fd_sc_hd__xor2_1
XU$$885 U$$885/A U$$929/B VGND VGND VPWR VPWR U$$885/X sky130_fd_sc_hd__xor2_1
XFILLER_44_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1035 U$$1446/A1 U$$1057/A2 U$$1448/A1 U$$1057/B2 VGND VGND VPWR VPWR U$$1036/A
+ sky130_fd_sc_hd__a22o_1
XU$$896 U$$896/A1 U$$938/A2 U$$896/B1 U$$938/B2 VGND VGND VPWR VPWR U$$897/A sky130_fd_sc_hd__a22o_1
XFILLER_31_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1046 U$$1046/A U$$968/B VGND VGND VPWR VPWR U$$1046/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1057 U$$98/A1 U$$1057/A2 U$$98/B1 U$$1057/B2 VGND VGND VPWR VPWR U$$1058/A sky130_fd_sc_hd__a22o_1
XU$$1068 U$$1068/A U$$962/A VGND VGND VPWR VPWR U$$1068/X sky130_fd_sc_hd__xor2_1
XFILLER_32_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1079 U$$2449/A1 U$$1093/A2 U$$1764/B1 U$$1093/B2 VGND VGND VPWR VPWR U$$1080/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_670 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_984 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_98_4 U$$3927/X U$$4060/X U$$4193/X VGND VGND VPWR VPWR dadda_fa_3_99_2/A
+ dadda_fa_3_98_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_171_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_41_0 U$$1552/X U$$1685/X U$$1818/X VGND VGND VPWR VPWR dadda_fa_3_42_0/B
+ dadda_fa_3_41_2/B sky130_fd_sc_hd__fa_1
XFILLER_39_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2270 U$$3366/A1 U$$2308/A2 U$$3366/B1 U$$2308/B2 VGND VGND VPWR VPWR U$$2271/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2281 U$$2281/A U$$2317/B VGND VGND VPWR VPWR U$$2281/X sky130_fd_sc_hd__xor2_1
XU$$2292 U$$2701/B1 U$$2316/A2 U$$2292/B1 U$$2316/B2 VGND VGND VPWR VPWR U$$2293/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1580 U$$1580/A U$$1620/B VGND VGND VPWR VPWR U$$1580/X sky130_fd_sc_hd__xor2_1
XU$$1591 U$$2550/A1 U$$1591/A2 U$$2415/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1592/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_70_2 dadda_fa_4_70_2/A dadda_fa_4_70_2/B dadda_fa_4_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_71_0/CIN dadda_fa_5_70_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_86_2 U$$2307/X U$$2440/X U$$2573/X VGND VGND VPWR VPWR dadda_fa_2_87_3/B
+ dadda_fa_2_86_5/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_63_1 dadda_fa_4_63_1/A dadda_fa_4_63_1/B dadda_fa_4_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/B dadda_fa_5_63_1/B sky130_fd_sc_hd__fa_1
XFILLER_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_79_1 U$$1495/X U$$1628/X U$$1761/X VGND VGND VPWR VPWR dadda_fa_2_80_0/CIN
+ dadda_fa_2_79_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_77_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_40_0 dadda_fa_7_40_0/A dadda_fa_7_40_0/B dadda_fa_7_40_0/CIN VGND VGND
+ VPWR VPWR _337_/D _208_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_56_0 dadda_fa_4_56_0/A dadda_fa_4_56_0/B dadda_fa_4_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/A dadda_fa_5_56_1/A sky130_fd_sc_hd__fa_1
XFILLER_58_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$210 final_adder.U$$210/A final_adder.U$$210/B VGND VGND VPWR VPWR
+ final_adder.U$$338/B sky130_fd_sc_hd__and2_1
XFILLER_57_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$221 final_adder.U$$220/B final_adder.U$$991/B1 final_adder.U$$221/B1
+ VGND VGND VPWR VPWR final_adder.U$$221/X sky130_fd_sc_hd__a21o_1
XTAP_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$232 final_adder.U$$232/A final_adder.U$$232/B VGND VGND VPWR VPWR
+ final_adder.U$$360/B sky130_fd_sc_hd__and2_1
XTAP_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$243 final_adder.U$$242/B final_adder.U$$243/A2 final_adder.U$$243/B1
+ VGND VGND VPWR VPWR final_adder.U$$243/X sky130_fd_sc_hd__a21o_1
XTAP_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$265 final_adder.U$$264/B final_adder.U$$139/X final_adder.U$$137/X
+ VGND VGND VPWR VPWR final_adder.U$$265/X sky130_fd_sc_hd__a21o_1
XTAP_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$104 U$$926/A1 U$$134/A2 U$$654/A1 U$$134/B2 VGND VGND VPWR VPWR U$$105/A sky130_fd_sc_hd__a22o_1
XFILLER_150_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$276 final_adder.U$$278/B final_adder.U$$276/B VGND VGND VPWR VPWR
+ final_adder.U$$402/B sky130_fd_sc_hd__and2_1
XU$$115 U$$115/A U$$127/B VGND VGND VPWR VPWR U$$115/X sky130_fd_sc_hd__xor2_1
XTAP_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater480 U$$3479/A2 VGND VGND VPWR VPWR U$$3453/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$287 final_adder.U$$286/B final_adder.U$$161/X final_adder.U$$159/X
+ VGND VGND VPWR VPWR final_adder.U$$287/X sky130_fd_sc_hd__a21o_1
Xrepeater491 U$$3416/A2 VGND VGND VPWR VPWR U$$3422/A2 sky130_fd_sc_hd__buf_6
XTAP_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$126 U$$674/A1 U$$134/A2 U$$950/A1 U$$134/B2 VGND VGND VPWR VPWR U$$127/A sky130_fd_sc_hd__a22o_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$298 final_adder.U$$300/B final_adder.U$$298/B VGND VGND VPWR VPWR
+ final_adder.U$$424/B sky130_fd_sc_hd__and2_1
XTAP_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$137 U$$3/A VGND VGND VPWR VPWR U$$137/Y sky130_fd_sc_hd__inv_1
XFILLER_72_334 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$148 U$$148/A U$$160/B VGND VGND VPWR VPWR U$$148/X sky130_fd_sc_hd__xor2_1
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$159 U$$22/A1 U$$165/A2 U$$24/A1 U$$165/B2 VGND VGND VPWR VPWR U$$160/A sky130_fd_sc_hd__a22o_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_392_ _401_/CLK _392_/D VGND VGND VPWR VPWR _392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1084 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1004 U$$4176/B1 VGND VGND VPWR VPWR U$$3902/B1 sky130_fd_sc_hd__buf_6
Xrepeater1015 input87/X VGND VGND VPWR VPWR U$$3846/B1 sky130_fd_sc_hd__buf_4
XFILLER_182_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_667 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1026 U$$3213/B1 VGND VGND VPWR VPWR U$$62/B1 sky130_fd_sc_hd__buf_6
XFILLER_114_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1037 input84/X VGND VGND VPWR VPWR U$$3211/B1 sky130_fd_sc_hd__buf_8
Xrepeater1048 input83/X VGND VGND VPWR VPWR U$$3485/A1 sky130_fd_sc_hd__buf_6
Xrepeater1059 U$$741/A1 VGND VGND VPWR VPWR U$$330/A1 sky130_fd_sc_hd__buf_6
XFILLER_181_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_426 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_74_0 dadda_fa_0_74_0/A U$$820/X U$$953/X VGND VGND VPWR VPWR dadda_fa_1_75_7/CIN
+ dadda_fa_1_74_8/B sky130_fd_sc_hd__fa_1
XFILLER_0_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput250 c[94] VGND VGND VPWR VPWR input250/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$660 U$$660/A1 U$$678/A2 U$$660/B1 U$$678/B2 VGND VGND VPWR VPWR U$$661/A sky130_fd_sc_hd__a22o_1
XU$$671 U$$671/A U$$685/A VGND VGND VPWR VPWR U$$671/X sky130_fd_sc_hd__xor2_1
XFILLER_56_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$682 U$$956/A1 U$$552/X U$$682/B1 U$$553/X VGND VGND VPWR VPWR U$$683/A sky130_fd_sc_hd__a22o_1
XU$$693 U$$967/A1 U$$711/A2 U$$969/A1 U$$711/B2 VGND VGND VPWR VPWR U$$694/A sky130_fd_sc_hd__a22o_1
XFILLER_189_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_80_1 dadda_fa_5_80_1/A dadda_fa_5_80_1/B dadda_fa_5_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_81_0/B dadda_fa_7_80_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_96_1 U$$2859/X U$$2992/X U$$3125/X VGND VGND VPWR VPWR dadda_fa_3_97_0/CIN
+ dadda_fa_3_96_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_73_0 dadda_fa_5_73_0/A dadda_fa_5_73_0/B dadda_fa_5_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_74_0/A dadda_fa_6_73_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1560 U$$4506/A1 VGND VGND VPWR VPWR U$$1764/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_154_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_89_0 U$$3377/X U$$3510/X U$$3643/X VGND VGND VPWR VPWR dadda_fa_3_90_0/B
+ dadda_fa_3_89_2/B sky130_fd_sc_hd__fa_1
Xrepeater1571 U$$3680/A1 VGND VGND VPWR VPWR U$$392/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_67_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1582 U$$2582/A1 VGND VGND VPWR VPWR U$$527/A1 sky130_fd_sc_hd__buf_4
Xrepeater1593 input113/X VGND VGND VPWR VPWR U$$3813/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_1_72_8 dadda_fa_1_72_8/A dadda_fa_1_72_8/B dadda_fa_1_72_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_73_3/A dadda_fa_3_72_0/A sky130_fd_sc_hd__fa_1
XFILLER_59_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_1188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_65_7 dadda_fa_1_65_7/A dadda_fa_1_65_7/B dadda_fa_1_65_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_2/CIN dadda_fa_2_65_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_802 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_6 U$$3980/X U$$4012/B input210/X VGND VGND VPWR VPWR dadda_fa_2_59_2/B
+ dadda_fa_2_58_5/B sky130_fd_sc_hd__fa_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_1_92_2 U$$2718/X U$$2851/X VGND VGND VPWR VPWR dadda_fa_2_93_5/B dadda_fa_3_92_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_88_0 dadda_fa_7_88_0/A dadda_fa_7_88_0/B dadda_fa_7_88_0/CIN VGND VGND
+ VPWR VPWR _385_/D _256_/D sky130_fd_sc_hd__fa_2
XFILLER_109_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_91_0 U$$1917/Y U$$2051/X U$$2184/X VGND VGND VPWR VPWR dadda_fa_2_92_4/B
+ dadda_fa_2_91_5/B sky130_fd_sc_hd__fa_1
XFILLER_159_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4408 U$$4408/A1 U$$4388/X U$$4408/B1 U$$4430/B2 VGND VGND VPWR VPWR U$$4409/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4419 U$$4419/A U$$4419/B VGND VGND VPWR VPWR U$$4419/X sky130_fd_sc_hd__xor2_1
XTAP_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3707 U$$3979/B1 U$$3793/A2 U$$832/A1 U$$3793/B2 VGND VGND VPWR VPWR U$$3708/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3718 U$$3718/A U$$3754/B VGND VGND VPWR VPWR U$$3718/X sky130_fd_sc_hd__xor2_1
XTAP_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3729 U$$4275/B1 U$$3773/A2 U$$4277/B1 U$$3773/B2 VGND VGND VPWR VPWR U$$3730/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_103_0 dadda_fa_6_103_0/A dadda_fa_6_103_0/B dadda_fa_6_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_104_0/B dadda_fa_7_103_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_23_3 U$$1516/X input172/X dadda_fa_3_23_3/CIN VGND VGND VPWR VPWR dadda_fa_4_24_1/B
+ dadda_fa_4_23_2/CIN sky130_fd_sc_hd__fa_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_375_ _377_/CLK _375_/D VGND VGND VPWR VPWR _375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_90_0 dadda_fa_6_90_0/A dadda_fa_6_90_0/B dadda_fa_6_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_91_0/B dadda_fa_7_90_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_10_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3568_1751 VGND VGND VPWR VPWR U$$3568_1751/HI U$$3568/A1 sky130_fd_sc_hd__conb_1
XFILLER_177_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_68_5 dadda_fa_2_68_5/A dadda_fa_2_68_5/B dadda_fa_2_68_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_69_2/A dadda_fa_4_68_0/A sky130_fd_sc_hd__fa_1
XFILLER_1_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1014 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$490 U$$490/A U$$492/B VGND VGND VPWR VPWR U$$490/X sky130_fd_sc_hd__xor2_1
XFILLER_211_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_954 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1390 U$$2454/B VGND VGND VPWR VPWR U$$2465/A sky130_fd_sc_hd__buf_6
XFILLER_120_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_70_5 U$$4270/X U$$4403/X input224/X VGND VGND VPWR VPWR dadda_fa_2_71_2/A
+ dadda_fa_2_70_5/A sky130_fd_sc_hd__fa_1
XFILLER_101_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_4 U$$3990/X U$$4123/X U$$4256/X VGND VGND VPWR VPWR dadda_fa_2_64_1/CIN
+ dadda_fa_2_63_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_56_3 U$$2380/X U$$2513/X U$$2646/X VGND VGND VPWR VPWR dadda_fa_2_57_1/B
+ dadda_fa_2_56_4/B sky130_fd_sc_hd__fa_1
XFILLER_132_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_33_2 dadda_fa_4_33_2/A dadda_fa_4_33_2/B dadda_fa_4_33_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_34_0/CIN dadda_fa_5_33_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_49_2 U$$903/X U$$1036/X U$$1169/X VGND VGND VPWR VPWR dadda_fa_2_50_1/B
+ dadda_fa_2_49_4/B sky130_fd_sc_hd__fa_1
XFILLER_131_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_26_1 dadda_fa_4_26_1/A dadda_fa_4_26_1/B dadda_fa_4_26_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/B dadda_fa_5_26_1/B sky130_fd_sc_hd__fa_1
XFILLER_199_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_0 U$$1109/X U$$1242/X input167/X VGND VGND VPWR VPWR dadda_fa_5_20_0/A
+ dadda_fa_5_19_1/A sky130_fd_sc_hd__fa_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_746 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_526 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2472_1733 VGND VGND VPWR VPWR U$$2472_1733/HI U$$2472/A1 sky130_fd_sc_hd__conb_1
XU$$4205 U$$4205/A U$$4227/B VGND VGND VPWR VPWR U$$4205/X sky130_fd_sc_hd__xor2_1
XU$$4216 U$$4490/A1 U$$4240/A2 U$$4492/A1 U$$4240/B2 VGND VGND VPWR VPWR U$$4217/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4227 U$$4227/A U$$4227/B VGND VGND VPWR VPWR U$$4227/X sky130_fd_sc_hd__xor2_1
XU$$4238 U$$4512/A1 U$$4238/A2 U$$4375/B1 U$$4238/B2 VGND VGND VPWR VPWR U$$4239/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3504 U$$3504/A U$$3504/B VGND VGND VPWR VPWR U$$3504/X sky130_fd_sc_hd__xor2_1
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4249 input60/X VGND VGND VPWR VPWR U$$4249/Y sky130_fd_sc_hd__inv_1
XU$$3515 U$$4335/B1 U$$3559/A2 U$$3517/A1 U$$3559/B2 VGND VGND VPWR VPWR U$$3516/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3526 U$$3526/A U$$3528/B VGND VGND VPWR VPWR U$$3526/X sky130_fd_sc_hd__xor2_1
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3537 input112/X U$$3559/A2 U$$3813/A1 U$$3559/B2 VGND VGND VPWR VPWR U$$3538/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3548 U$$3548/A U$$3550/B VGND VGND VPWR VPWR U$$3548/X sky130_fd_sc_hd__xor2_1
XU$$2803 U$$2803/A U$$2825/B VGND VGND VPWR VPWR U$$2803/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3559 input124/X U$$3559/A2 U$$3559/B1 U$$3559/B2 VGND VGND VPWR VPWR U$$3560/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2814 U$$2951/A1 U$$2828/A2 U$$2951/B1 U$$2828/B2 VGND VGND VPWR VPWR U$$2815/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2825 U$$2825/A U$$2825/B VGND VGND VPWR VPWR U$$2825/X sky130_fd_sc_hd__xor2_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2836 U$$3108/B1 U$$2844/A2 U$$2975/A1 U$$2844/B2 VGND VGND VPWR VPWR U$$2837/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_3_21_0 U$$49/X U$$182/X U$$315/X VGND VGND VPWR VPWR dadda_fa_4_22_0/B dadda_fa_4_21_1/CIN
+ sky130_fd_sc_hd__fa_1
XU$$2847 U$$2847/A U$$2876/A VGND VGND VPWR VPWR U$$2847/X sky130_fd_sc_hd__xor2_1
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2858 U$$3680/A1 U$$2858/A2 U$$118/B1 U$$2858/B2 VGND VGND VPWR VPWR U$$2859/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 U$$2828/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2869 U$$2869/A U$$2869/B VGND VGND VPWR VPWR U$$2869/X sky130_fd_sc_hd__xor2_1
XANTENNA_152 U$$3227/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_196 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1064 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1026 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_358_ _358_/CLK _358_/D VGND VGND VPWR VPWR _358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_289_ _419_/CLK _289_/D VGND VGND VPWR VPWR _289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_80_4 dadda_fa_2_80_4/A dadda_fa_2_80_4/B dadda_fa_2_80_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_1/CIN dadda_fa_3_80_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_73_3 dadda_fa_2_73_3/A dadda_fa_2_73_3/B dadda_fa_2_73_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/B dadda_fa_3_73_3/B sky130_fd_sc_hd__fa_1
XFILLER_29_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_66_2 dadda_fa_2_66_2/A dadda_fa_2_66_2/B dadda_fa_2_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/A dadda_fa_3_66_3/A sky130_fd_sc_hd__fa_2
XFILLER_68_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$809 final_adder.U$$776/A final_adder.U$$729/X final_adder.U$$697/X
+ VGND VGND VPWR VPWR final_adder.U$$809/X sky130_fd_sc_hd__a21o_1
XFILLER_57_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_43_1 dadda_fa_5_43_1/A dadda_fa_5_43_1/B dadda_fa_5_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_44_0/B dadda_fa_7_43_0/A sky130_fd_sc_hd__fa_2
XFILLER_84_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_727 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_59_1 dadda_fa_2_59_1/A dadda_fa_2_59_1/B dadda_fa_2_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_0/CIN dadda_fa_3_59_2/CIN sky130_fd_sc_hd__fa_1
Xinput3 a[11] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_4
Xdadda_fa_5_36_0 dadda_fa_5_36_0/A dadda_fa_5_36_0/B dadda_fa_5_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_37_0/A dadda_fa_6_36_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_37_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4495_1824 VGND VGND VPWR VPWR U$$4495_1824/HI U$$4495/B sky130_fd_sc_hd__conb_1
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_110_0 dadda_fa_5_110_0/A dadda_fa_5_110_0/B dadda_fa_5_110_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_111_0/A dadda_fa_6_110_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1 _297_/Q _169_/Q VGND VGND VPWR VPWR final_adder.U$$255/B1 final_adder.U$$1/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_152_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_581 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput340 output340/A VGND VGND VPWR VPWR o[5] sky130_fd_sc_hd__buf_2
XFILLER_134_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput351 output351/A VGND VGND VPWR VPWR o[6] sky130_fd_sc_hd__buf_2
Xoutput362 output362/A VGND VGND VPWR VPWR o[7] sky130_fd_sc_hd__buf_2
XFILLER_105_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput373 output373/A VGND VGND VPWR VPWR o[8] sky130_fd_sc_hd__buf_2
XFILLER_121_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_275 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput384 output384/A VGND VGND VPWR VPWR o[9] sky130_fd_sc_hd__buf_2
XFILLER_43_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_61_1 U$$2390/X U$$2523/X U$$2656/X VGND VGND VPWR VPWR dadda_fa_2_62_0/CIN
+ dadda_fa_2_61_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_54_0 U$$780/X U$$913/X U$$1046/X VGND VGND VPWR VPWR dadda_fa_2_55_0/B
+ dadda_fa_2_54_3/B sky130_fd_sc_hd__fa_1
XFILLER_28_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1409 U$$1409/A U$$1423/B VGND VGND VPWR VPWR U$$1409/X sky130_fd_sc_hd__xor2_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1015 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_212_ _219_/CLK _212_/D VGND VGND VPWR VPWR _212_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_204_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_90_3 dadda_fa_3_90_3/A dadda_fa_3_90_3/B dadda_fa_3_90_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_91_1/B dadda_fa_4_90_2/CIN sky130_fd_sc_hd__fa_2
XFILLER_87_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_83_2 dadda_fa_3_83_2/A dadda_fa_3_83_2/B dadda_fa_3_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_1/A dadda_fa_4_83_2/B sky130_fd_sc_hd__fa_1
XFILLER_139_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_76_1 dadda_fa_3_76_1/A dadda_fa_3_76_1/B dadda_fa_3_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_0/CIN dadda_fa_4_76_2/A sky130_fd_sc_hd__fa_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_53_0 dadda_fa_6_53_0/A dadda_fa_6_53_0/B dadda_fa_6_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_54_0/B dadda_fa_7_53_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_69_0 dadda_fa_3_69_0/A dadda_fa_3_69_0/B dadda_fa_3_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_0/B dadda_fa_4_69_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_111_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4002 U$$4002/A U$$4036/B VGND VGND VPWR VPWR U$$4002/X sky130_fd_sc_hd__xor2_1
XU$$4013 input72/X U$$4079/A2 U$$4013/B1 U$$4079/B2 VGND VGND VPWR VPWR U$$4014/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4024 U$$4024/A U$$4109/A VGND VGND VPWR VPWR U$$4024/X sky130_fd_sc_hd__xor2_1
XU$$4035 U$$4309/A1 U$$4035/A2 U$$4309/B1 U$$4035/B2 VGND VGND VPWR VPWR U$$4036/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4046 U$$4046/A U$$4100/B VGND VGND VPWR VPWR U$$4046/X sky130_fd_sc_hd__xor2_1
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3301 U$$3301/A U$$3321/B VGND VGND VPWR VPWR U$$3301/X sky130_fd_sc_hd__xor2_1
XU$$4057 U$$4466/B1 U$$4077/A2 U$$4333/A1 U$$4077/B2 VGND VGND VPWR VPWR U$$4058/A
+ sky130_fd_sc_hd__a22o_1
XU$$3312 U$$4408/A1 U$$3348/A2 input128/X U$$3394/B2 VGND VGND VPWR VPWR U$$3313/A
+ sky130_fd_sc_hd__a22o_1
XU$$4068 U$$4068/A U$$4078/B VGND VGND VPWR VPWR U$$4068/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_112_2 dadda_fa_4_112_2/A dadda_fa_4_112_2/B dadda_ha_3_112_2/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_113_0/CIN dadda_fa_5_112_1/CIN sky130_fd_sc_hd__fa_1
XU$$3323 U$$3323/A U$$3349/B VGND VGND VPWR VPWR U$$3323/X sky130_fd_sc_hd__xor2_1
XU$$3334 U$$4430/A1 U$$3374/A2 U$$4432/A1 U$$3374/B2 VGND VGND VPWR VPWR U$$3335/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4079 U$$517/A1 U$$4079/A2 U$$517/B1 U$$4079/B2 VGND VGND VPWR VPWR U$$4080/A sky130_fd_sc_hd__a22o_1
XFILLER_206_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2600 U$$3148/A1 U$$2600/A2 U$$2600/B1 U$$2600/B2 VGND VGND VPWR VPWR U$$2601/A
+ sky130_fd_sc_hd__a22o_1
XU$$3345 U$$3345/A U$$3425/A VGND VGND VPWR VPWR U$$3345/X sky130_fd_sc_hd__xor2_1
XFILLER_18_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2611 U$$3159/A1 U$$2625/A2 U$$3296/B1 U$$2625/B2 VGND VGND VPWR VPWR U$$2612/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3356 U$$3356/A1 U$$3388/A2 U$$4178/B1 U$$3378/B2 VGND VGND VPWR VPWR U$$3357/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_105_1 dadda_fa_4_105_1/A dadda_fa_4_105_1/B dadda_fa_4_105_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/B dadda_fa_5_105_1/B sky130_fd_sc_hd__fa_1
XU$$3367 U$$3367/A U$$3377/B VGND VGND VPWR VPWR U$$3367/X sky130_fd_sc_hd__xor2_1
XU$$2622 U$$2622/A U$$2624/B VGND VGND VPWR VPWR U$$2622/X sky130_fd_sc_hd__xor2_1
XFILLER_62_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2633 U$$578/A1 U$$2653/A2 U$$3183/A1 U$$2653/B2 VGND VGND VPWR VPWR U$$2634/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3378 U$$3378/A1 U$$3378/A2 U$$3517/A1 U$$3378/B2 VGND VGND VPWR VPWR U$$3379/A
+ sky130_fd_sc_hd__a22o_1
XU$$2644 U$$2644/A U$$2650/B VGND VGND VPWR VPWR U$$2644/X sky130_fd_sc_hd__xor2_1
XFILLER_62_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3389 U$$3389/A U$$3389/B VGND VGND VPWR VPWR U$$3389/X sky130_fd_sc_hd__xor2_1
XU$$1910 U$$1910/A U$$1912/B VGND VGND VPWR VPWR U$$1910/X sky130_fd_sc_hd__xor2_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2655 U$$463/A1 U$$2683/A2 U$$874/B1 U$$2683/B2 VGND VGND VPWR VPWR U$$2656/A sky130_fd_sc_hd__a22o_1
XU$$2666 U$$2666/A U$$2710/B VGND VGND VPWR VPWR U$$2666/X sky130_fd_sc_hd__xor2_1
XFILLER_34_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1921 U$$2047/B U$$1921/B VGND VGND VPWR VPWR U$$1921/X sky130_fd_sc_hd__and2_1
XFILLER_92_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2677 U$$3088/A1 U$$2691/A2 U$$3499/B1 U$$2691/B2 VGND VGND VPWR VPWR U$$2678/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1932 U$$2069/A1 U$$1970/A2 U$$1932/B1 U$$1970/B2 VGND VGND VPWR VPWR U$$1933/A
+ sky130_fd_sc_hd__a22o_1
XU$$2688 U$$2688/A U$$2739/A VGND VGND VPWR VPWR U$$2688/X sky130_fd_sc_hd__xor2_1
XU$$1943 U$$1943/A U$$1991/B VGND VGND VPWR VPWR U$$1943/X sky130_fd_sc_hd__xor2_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1954 U$$4009/A1 U$$1960/A2 U$$860/A1 U$$1960/B2 VGND VGND VPWR VPWR U$$1955/A
+ sky130_fd_sc_hd__a22o_1
XU$$2699 U$$3245/B1 U$$2711/A2 U$$3112/A1 U$$2711/B2 VGND VGND VPWR VPWR U$$2700/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1965 U$$1965/A U$$1991/B VGND VGND VPWR VPWR U$$1965/X sky130_fd_sc_hd__xor2_1
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1976 U$$3618/B1 U$$2016/A2 U$$2113/B1 U$$2016/B2 VGND VGND VPWR VPWR U$$1977/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_126_0 dadda_fa_7_126_0/A dadda_fa_7_126_0/B dadda_fa_7_126_0/CIN VGND
+ VGND VPWR VPWR _423_/D _294_/D sky130_fd_sc_hd__fa_1
XU$$1987 U$$1987/A U$$2017/B VGND VGND VPWR VPWR U$$1987/X sky130_fd_sc_hd__xor2_1
XFILLER_109_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1998 U$$3366/B1 U$$2040/A2 U$$2409/B1 U$$2040/B2 VGND VGND VPWR VPWR U$$1999/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_71_0 dadda_fa_2_71_0/A dadda_fa_2_71_0/B dadda_fa_2_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_0/B dadda_fa_3_71_2/B sky130_fd_sc_hd__fa_1
XFILLER_102_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_100_0_1860 VGND VGND VPWR VPWR dadda_fa_2_100_0/A dadda_fa_2_100_0_1860/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_29_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$606 final_adder.U$$614/B final_adder.U$$606/B VGND VGND VPWR VPWR
+ final_adder.U$$710/A sky130_fd_sc_hd__and2_1
Xrepeater810 U$$2326/B2 VGND VGND VPWR VPWR U$$2284/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$617 final_adder.U$$616/B final_adder.U$$501/X final_adder.U$$493/X
+ VGND VGND VPWR VPWR final_adder.U$$617/X sky130_fd_sc_hd__a21o_1
Xrepeater821 U$$2060/X VGND VGND VPWR VPWR U$$2169/B2 sky130_fd_sc_hd__buf_6
XFILLER_84_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$628 final_adder.U$$644/B final_adder.U$$628/B VGND VGND VPWR VPWR
+ final_adder.U$$740/B sky130_fd_sc_hd__and2_1
XFILLER_57_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater832 U$$1879/B2 VGND VGND VPWR VPWR U$$1831/B2 sky130_fd_sc_hd__buf_8
Xfinal_adder.U$$639 final_adder.U$$638/B final_adder.U$$535/X final_adder.U$$519/X
+ VGND VGND VPWR VPWR final_adder.U$$639/X sky130_fd_sc_hd__a21o_1
Xrepeater843 U$$1746/B2 VGND VGND VPWR VPWR U$$1750/B2 sky130_fd_sc_hd__buf_4
XFILLER_42_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater854 U$$1512/X VGND VGND VPWR VPWR U$$1637/B2 sky130_fd_sc_hd__buf_6
Xrepeater865 U$$1422/B2 VGND VGND VPWR VPWR U$$1404/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_99_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater876 U$$1291/B2 VGND VGND VPWR VPWR U$$1281/B2 sky130_fd_sc_hd__clkbuf_4
Xrepeater887 U$$94/B2 VGND VGND VPWR VPWR U$$98/B2 sky130_fd_sc_hd__buf_6
Xrepeater898 U$$4498/B2 VGND VGND VPWR VPWR U$$4476/B2 sky130_fd_sc_hd__buf_4
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$50 U$$50/A1 U$$50/A2 U$$52/A1 U$$50/B2 VGND VGND VPWR VPWR U$$51/A sky130_fd_sc_hd__a22o_1
XU$$61 U$$61/A U$$85/B VGND VGND VPWR VPWR U$$61/X sky130_fd_sc_hd__xor2_1
XFILLER_112_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$72 U$$72/A1 U$$80/A2 U$$74/A1 U$$80/B2 VGND VGND VPWR VPWR U$$73/A sky130_fd_sc_hd__a22o_1
XU$$83 U$$83/A U$$85/B VGND VGND VPWR VPWR U$$83/X sky130_fd_sc_hd__xor2_1
XFILLER_52_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$94 U$$94/A1 U$$94/A2 U$$96/A1 U$$94/B2 VGND VGND VPWR VPWR U$$95/A sky130_fd_sc_hd__a22o_1
XU$$3890 input80/X U$$3840/X U$$4029/A1 U$$3841/X VGND VGND VPWR VPWR U$$3891/A sky130_fd_sc_hd__a22o_1
XFILLER_13_808 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_30 _339_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_63 _342_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_74 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_4_93_1 dadda_fa_4_93_1/A dadda_fa_4_93_1/B dadda_fa_4_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/B dadda_fa_5_93_1/B sky130_fd_sc_hd__fa_1
XFILLER_10_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_88_0_1856 VGND VGND VPWR VPWR dadda_fa_1_88_0/A dadda_fa_1_88_0_1856/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_192_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_70_0 dadda_fa_7_70_0/A dadda_fa_7_70_0/B dadda_fa_7_70_0/CIN VGND VGND
+ VPWR VPWR _367_/D _238_/D sky130_fd_sc_hd__fa_1
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_86_0 dadda_fa_4_86_0/A dadda_fa_4_86_0/B dadda_fa_4_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/A dadda_fa_5_86_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_107_3 input137/X dadda_fa_3_107_3/B dadda_fa_3_107_3/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_108_1/B dadda_fa_4_107_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1063 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1206 U$$932/A1 U$$1100/X U$$932/B1 U$$1101/X VGND VGND VPWR VPWR U$$1207/A sky130_fd_sc_hd__a22o_1
XFILLER_71_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1217 U$$1217/A U$$1223/B VGND VGND VPWR VPWR U$$1217/X sky130_fd_sc_hd__xor2_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1228 U$$2324/A1 U$$1230/A2 U$$1504/A1 U$$1230/B2 VGND VGND VPWR VPWR U$$1229/A
+ sky130_fd_sc_hd__a22o_1
XU$$1239 U$$1239/A1 U$$1311/A2 U$$1515/A1 U$$1271/B2 VGND VGND VPWR VPWR U$$1240/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1011 final_adder.U$$240/A final_adder.U$$621/X final_adder.U$$241/A2
+ VGND VGND VPWR VPWR final_adder.U$$1039/B sky130_fd_sc_hd__a21o_1
XFILLER_141_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1033 final_adder.U$$9/SUM final_adder.U$$1033/B VGND VGND VPWR VPWR
+ output384/A sky130_fd_sc_hd__xor2_1
XFILLER_89_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1044 final_adder.U$$234/A final_adder.U$$735/X VGND VGND VPWR VPWR
+ output297/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1055 final_adder.U$$224/B final_adder.U$$995/X VGND VGND VPWR VPWR
+ output309/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1066 final_adder.U$$212/A final_adder.U$$825/X VGND VGND VPWR VPWR
+ output321/A sky130_fd_sc_hd__xor2_1
XFILLER_7_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1077 final_adder.U$$202/B final_adder.U$$973/X VGND VGND VPWR VPWR
+ output333/A sky130_fd_sc_hd__xor2_1
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1088 final_adder.U$$190/A final_adder.U$$803/X VGND VGND VPWR VPWR
+ output345/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1099 final_adder.U$$180/B final_adder.U$$951/X VGND VGND VPWR VPWR
+ output357/A sky130_fd_sc_hd__xor2_1
XFILLER_139_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1086 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_50_5 dadda_fa_2_50_5/A dadda_fa_2_50_5/B dadda_fa_2_50_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_51_2/A dadda_fa_4_50_0/A sky130_fd_sc_hd__fa_1
XFILLER_4_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_43_4 dadda_fa_2_43_4/A dadda_fa_2_43_4/B dadda_fa_2_43_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_1/CIN dadda_fa_3_43_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3120 U$$517/A1 U$$3132/A2 U$$517/B1 U$$3132/B2 VGND VGND VPWR VPWR U$$3121/A sky130_fd_sc_hd__a22o_1
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3131 U$$3131/A U$$3133/B VGND VGND VPWR VPWR U$$3131/X sky130_fd_sc_hd__xor2_1
XFILLER_4_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3142 input121/X U$$3148/A2 U$$3281/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3143/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_6_2_0 U$$11/X U$$144/X VGND VGND VPWR VPWR dadda_fa_7_3_0/B dadda_ha_6_2_0/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_59_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3153 U$$3288/A VGND VGND VPWR VPWR U$$3153/Y sky130_fd_sc_hd__inv_1
XFILLER_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_36_3 U$$1941/X U$$2074/X U$$2207/X VGND VGND VPWR VPWR dadda_fa_3_37_1/B
+ dadda_fa_3_36_3/B sky130_fd_sc_hd__fa_1
XFILLER_81_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3164 U$$3164/A U$$3188/B VGND VGND VPWR VPWR U$$3164/X sky130_fd_sc_hd__xor2_1
XFILLER_207_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3175 input127/X U$$3263/A2 U$$3451/A1 U$$3263/B2 VGND VGND VPWR VPWR U$$3176/A
+ sky130_fd_sc_hd__a22o_1
XU$$2430 U$$2430/A U$$2454/B VGND VGND VPWR VPWR U$$2430/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2441 U$$934/A1 U$$2333/X U$$936/A1 U$$2334/X VGND VGND VPWR VPWR U$$2442/A sky130_fd_sc_hd__a22o_1
XU$$3186 U$$3186/A U$$3188/B VGND VGND VPWR VPWR U$$3186/X sky130_fd_sc_hd__xor2_1
XU$$2452 U$$2452/A U$$2454/B VGND VGND VPWR VPWR U$$2452/X sky130_fd_sc_hd__xor2_1
XU$$3197 U$$4430/A1 U$$3241/A2 U$$4432/A1 U$$3241/B2 VGND VGND VPWR VPWR U$$3198/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2463 U$$3148/A1 U$$2463/A2 U$$2463/B1 U$$2463/B2 VGND VGND VPWR VPWR U$$2464/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_29_2 U$$863/X U$$996/X U$$1129/X VGND VGND VPWR VPWR dadda_fa_3_30_2/A
+ dadda_fa_3_29_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2474 U$$2609/B1 U$$2524/A2 U$$3296/B1 U$$2524/B2 VGND VGND VPWR VPWR U$$2475/A
+ sky130_fd_sc_hd__a22o_1
XU$$2485 U$$2485/A U$$2491/B VGND VGND VPWR VPWR U$$2485/X sky130_fd_sc_hd__xor2_1
XU$$1740 U$$96/A1 U$$1746/A2 U$$2016/A1 U$$1746/B2 VGND VGND VPWR VPWR U$$1741/A sky130_fd_sc_hd__a22o_1
XFILLER_210_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1751 U$$1751/A U$$1751/B VGND VGND VPWR VPWR U$$1751/X sky130_fd_sc_hd__xor2_1
XU$$2496 U$$989/A1 U$$2542/A2 U$$3183/A1 U$$2542/B2 VGND VGND VPWR VPWR U$$2497/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1762 U$$527/B1 U$$1764/A2 U$$2312/A1 U$$1764/B2 VGND VGND VPWR VPWR U$$1763/A
+ sky130_fd_sc_hd__a22o_1
XU$$1773 U$$1773/A U$$1779/B VGND VGND VPWR VPWR U$$1773/X sky130_fd_sc_hd__xor2_1
XU$$1784 input20/X U$$1784/B VGND VGND VPWR VPWR U$$1784/X sky130_fd_sc_hd__and2_1
XFILLER_210_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1795 U$$2343/A1 U$$1819/A2 U$$1932/B1 U$$1819/B2 VGND VGND VPWR VPWR U$$1796/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_0_76_0_1851 VGND VGND VPWR VPWR dadda_fa_0_76_0/A dadda_fa_0_76_0_1851/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_162_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput50 a[54] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_1
Xinput61 a[6] VGND VGND VPWR VPWR U$$412/A sky130_fd_sc_hd__buf_2
Xinput72 b[16] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__buf_8
XFILLER_174_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput83 b[26] VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_8
Xinput94 b[36] VGND VGND VPWR VPWR input94/X sky130_fd_sc_hd__buf_6
XFILLER_157_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$403 final_adder.U$$402/B final_adder.U$$281/X final_adder.U$$277/X
+ VGND VGND VPWR VPWR final_adder.U$$403/X sky130_fd_sc_hd__a21o_1
XTAP_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$414 final_adder.U$$418/B final_adder.U$$414/B VGND VGND VPWR VPWR
+ final_adder.U$$538/B sky130_fd_sc_hd__and2_1
XFILLER_112_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$425 final_adder.U$$424/B final_adder.U$$303/X final_adder.U$$299/X
+ VGND VGND VPWR VPWR final_adder.U$$425/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$436 final_adder.U$$440/B final_adder.U$$436/B VGND VGND VPWR VPWR
+ final_adder.U$$560/B sky130_fd_sc_hd__and2_1
XTAP_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater640 U$$1083/B2 VGND VGND VPWR VPWR U$$993/B2 sky130_fd_sc_hd__buf_4
XFILLER_111_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$447 final_adder.U$$446/B final_adder.U$$325/X final_adder.U$$321/X
+ VGND VGND VPWR VPWR final_adder.U$$447/X sky130_fd_sc_hd__a21o_1
XTAP_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater651 U$$950/B2 VGND VGND VPWR VPWR U$$906/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$458 final_adder.U$$462/B final_adder.U$$458/B VGND VGND VPWR VPWR
+ final_adder.U$$582/B sky130_fd_sc_hd__and2_1
XTAP_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater662 U$$624/B2 VGND VGND VPWR VPWR U$$616/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$469 final_adder.U$$468/B final_adder.U$$347/X final_adder.U$$343/X
+ VGND VGND VPWR VPWR final_adder.U$$469/X sky130_fd_sc_hd__a21o_1
XU$$308 U$$34/A1 U$$316/A2 U$$36/A1 U$$316/B2 VGND VGND VPWR VPWR U$$309/A sky130_fd_sc_hd__a22o_1
XFILLER_57_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater673 U$$4369/B2 VGND VGND VPWR VPWR U$$4327/B2 sky130_fd_sc_hd__buf_4
Xrepeater684 U$$416/X VGND VGND VPWR VPWR U$$527/B2 sky130_fd_sc_hd__buf_6
XU$$319 U$$319/A U$$343/B VGND VGND VPWR VPWR U$$319/X sky130_fd_sc_hd__xor2_1
Xrepeater695 U$$4043/B2 VGND VGND VPWR VPWR U$$4035/B2 sky130_fd_sc_hd__buf_6
XFILLER_44_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_446 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1002 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1208 U$$684/A VGND VGND VPWR VPWR U$$637/B sky130_fd_sc_hd__buf_8
Xdadda_fa_3_112_1 U$$3689/X U$$3822/X U$$3955/X VGND VGND VPWR VPWR dadda_fa_4_113_1/CIN
+ dadda_fa_4_112_2/B sky130_fd_sc_hd__fa_1
Xrepeater1219 U$$528/B VGND VGND VPWR VPWR U$$516/B sky130_fd_sc_hd__buf_6
XFILLER_5_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_359 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_105_0 U$$3675/X U$$3808/X U$$3941/X VGND VGND VPWR VPWR dadda_fa_4_106_0/B
+ dadda_fa_4_105_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_134_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_53_3 dadda_fa_3_53_3/A dadda_fa_3_53_3/B dadda_fa_3_53_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_54_1/B dadda_fa_4_53_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_75_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_69_3 U$$1608/X U$$1741/X U$$1874/X VGND VGND VPWR VPWR dadda_fa_1_70_7/A
+ dadda_fa_1_69_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_209_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_46_2 dadda_fa_3_46_2/A dadda_fa_3_46_2/B dadda_fa_3_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_1/A dadda_fa_4_46_2/B sky130_fd_sc_hd__fa_1
XTAP_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$981 final_adder.U$$210/A final_adder.U$$823/X final_adder.U$$981/B1
+ VGND VGND VPWR VPWR final_adder.U$$981/X sky130_fd_sc_hd__a21o_1
XFILLER_180_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_39_1 dadda_fa_3_39_1/A dadda_fa_3_39_1/B dadda_fa_3_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_0/CIN dadda_fa_4_39_2/A sky130_fd_sc_hd__fa_1
XFILLER_90_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$820 U$$820/A U$$821/A VGND VGND VPWR VPWR U$$820/X sky130_fd_sc_hd__xor2_1
XU$$831 U$$831/A U$$847/B VGND VGND VPWR VPWR U$$831/X sky130_fd_sc_hd__xor2_1
XU$$842 U$$979/A1 U$$906/A2 U$$842/B1 U$$906/B2 VGND VGND VPWR VPWR U$$843/A sky130_fd_sc_hd__a22o_1
XFILLER_169_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_16_0 dadda_fa_6_16_0/A dadda_fa_6_16_0/B dadda_fa_6_16_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_17_0/B dadda_fa_7_16_0/CIN sky130_fd_sc_hd__fa_1
XU$$853 U$$853/A U$$877/B VGND VGND VPWR VPWR U$$853/X sky130_fd_sc_hd__xor2_1
XFILLER_204_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1003 U$$866/A1 U$$999/A2 U$$46/A1 U$$999/B2 VGND VGND VPWR VPWR U$$1004/A sky130_fd_sc_hd__a22o_1
XFILLER_44_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$864 U$$864/A1 U$$882/A2 U$$864/B1 U$$882/B2 VGND VGND VPWR VPWR U$$865/A sky130_fd_sc_hd__a22o_1
XFILLER_204_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1014 U$$1014/A U$$998/B VGND VGND VPWR VPWR U$$1014/X sky130_fd_sc_hd__xor2_1
XU$$875 U$$875/A U$$951/B VGND VGND VPWR VPWR U$$875/X sky130_fd_sc_hd__xor2_1
XFILLER_189_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$886 U$$62/B1 U$$892/A2 U$$888/A1 U$$892/B2 VGND VGND VPWR VPWR U$$887/A sky130_fd_sc_hd__a22o_1
XU$$1025 U$$888/A1 U$$993/A2 U$$890/A1 U$$993/B2 VGND VGND VPWR VPWR U$$1026/A sky130_fd_sc_hd__a22o_1
XFILLER_204_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$897 U$$897/A U$$945/B VGND VGND VPWR VPWR U$$897/X sky130_fd_sc_hd__xor2_1
XFILLER_44_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1036 U$$1036/A U$$980/B VGND VGND VPWR VPWR U$$1036/X sky130_fd_sc_hd__xor2_1
XFILLER_189_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1047 U$$910/A1 U$$965/A2 U$$912/A1 U$$965/B2 VGND VGND VPWR VPWR U$$1048/A sky130_fd_sc_hd__a22o_1
XFILLER_73_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1058 U$$1058/A U$$1084/B VGND VGND VPWR VPWR U$$1058/X sky130_fd_sc_hd__xor2_1
XFILLER_73_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1069 U$$2711/B1 U$$963/X U$$934/A1 U$$964/X VGND VGND VPWR VPWR U$$1070/A sky130_fd_sc_hd__a22o_1
XFILLER_148_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_446 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_41_1 U$$1951/X U$$2084/X U$$2217/X VGND VGND VPWR VPWR dadda_fa_3_42_0/CIN
+ dadda_fa_3_41_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_34_0 U$$341/X U$$474/X U$$607/X VGND VGND VPWR VPWR dadda_fa_3_35_0/B
+ dadda_fa_3_34_2/B sky130_fd_sc_hd__fa_1
XFILLER_207_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2260 U$$3356/A1 U$$2308/A2 U$$2808/B1 U$$2308/B2 VGND VGND VPWR VPWR U$$2261/A
+ sky130_fd_sc_hd__a22o_1
XU$$2271 U$$2271/A U$$2309/B VGND VGND VPWR VPWR U$$2271/X sky130_fd_sc_hd__xor2_1
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2282 U$$2282/A1 U$$2302/A2 U$$366/A1 U$$2302/B2 VGND VGND VPWR VPWR U$$2283/A
+ sky130_fd_sc_hd__a22o_1
XU$$2293 U$$2293/A U$$2317/B VGND VGND VPWR VPWR U$$2293/X sky130_fd_sc_hd__xor2_1
XFILLER_210_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1570 U$$1570/A U$$1574/B VGND VGND VPWR VPWR U$$1570/X sky130_fd_sc_hd__xor2_1
XU$$1581 U$$2951/A1 U$$1621/A2 U$$2951/B1 U$$1621/B2 VGND VGND VPWR VPWR U$$1582/A
+ sky130_fd_sc_hd__a22o_1
XU$$1592 U$$1592/A U$$1592/B VGND VGND VPWR VPWR U$$1592/X sky130_fd_sc_hd__xor2_1
XFILLER_148_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_86_3 U$$2706/X U$$2839/X U$$2972/X VGND VGND VPWR VPWR dadda_fa_2_87_3/CIN
+ dadda_fa_2_86_5/B sky130_fd_sc_hd__fa_1
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_63_2 dadda_fa_4_63_2/A dadda_fa_4_63_2/B dadda_fa_4_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_64_0/CIN dadda_fa_5_63_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_79_2 U$$1894/X U$$2027/X U$$2160/X VGND VGND VPWR VPWR dadda_fa_2_80_1/A
+ dadda_fa_2_79_4/A sky130_fd_sc_hd__fa_1
XFILLER_103_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_56_1 dadda_fa_4_56_1/A dadda_fa_4_56_1/B dadda_fa_4_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/B dadda_fa_5_56_1/B sky130_fd_sc_hd__fa_1
XTAP_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$200 final_adder.U$$200/A final_adder.U$$200/B VGND VGND VPWR VPWR
+ final_adder.U$$328/B sky130_fd_sc_hd__and2_1
XFILLER_170_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$211 final_adder.U$$210/B final_adder.U$$981/B1 final_adder.U$$211/B1
+ VGND VGND VPWR VPWR final_adder.U$$211/X sky130_fd_sc_hd__a21o_1
XTAP_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_33_0 dadda_fa_7_33_0/A dadda_fa_7_33_0/B dadda_fa_7_33_0/CIN VGND VGND
+ VPWR VPWR _330_/D _201_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$222 final_adder.U$$222/A final_adder.U$$222/B VGND VGND VPWR VPWR
+ final_adder.U$$350/B sky130_fd_sc_hd__and2_1
XTAP_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_49_0 dadda_fa_4_49_0/A dadda_fa_4_49_0/B dadda_fa_4_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/A dadda_fa_5_49_1/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$233 final_adder.U$$232/B final_adder.U$$233/A2 final_adder.U$$233/B1
+ VGND VGND VPWR VPWR final_adder.U$$233/X sky130_fd_sc_hd__a21o_1
XTAP_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$244 final_adder.U$$244/A final_adder.U$$244/B VGND VGND VPWR VPWR
+ final_adder.U$$372/B sky130_fd_sc_hd__and2_1
XTAP_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$255 final_adder.U$$1/SUM final_adder.U$$255/A2 final_adder.U$$255/B1
+ VGND VGND VPWR VPWR final_adder.U$$255/X sky130_fd_sc_hd__a21o_2
XTAP_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$266 final_adder.U$$268/B final_adder.U$$266/B VGND VGND VPWR VPWR
+ final_adder.U$$392/B sky130_fd_sc_hd__and2_1
XTAP_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater470 U$$3703/X VGND VGND VPWR VPWR U$$3777/A2 sky130_fd_sc_hd__buf_6
XU$$105 U$$105/A U$$111/B VGND VGND VPWR VPWR U$$105/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$277 final_adder.U$$276/B final_adder.U$$151/X final_adder.U$$149/X
+ VGND VGND VPWR VPWR final_adder.U$$277/X sky130_fd_sc_hd__a21o_1
XU$$116 U$$116/A1 U$$122/A2 U$$392/A1 U$$122/B2 VGND VGND VPWR VPWR U$$117/A sky130_fd_sc_hd__a22o_1
XTAP_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater481 U$$3429/X VGND VGND VPWR VPWR U$$3479/A2 sky130_fd_sc_hd__buf_6
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$288 final_adder.U$$290/B final_adder.U$$288/B VGND VGND VPWR VPWR
+ final_adder.U$$414/B sky130_fd_sc_hd__and2_1
XTAP_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$127 U$$127/A U$$127/B VGND VGND VPWR VPWR U$$127/X sky130_fd_sc_hd__xor2_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater492 U$$3388/A2 VGND VGND VPWR VPWR U$$3416/A2 sky130_fd_sc_hd__buf_6
XFILLER_84_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$299 final_adder.U$$298/B final_adder.U$$173/X final_adder.U$$171/X
+ VGND VGND VPWR VPWR final_adder.U$$299/X sky130_fd_sc_hd__a21o_1
XU$$138 U$$138/A VGND VGND VPWR VPWR U$$140/B sky130_fd_sc_hd__inv_1
XU$$149 U$$12/A1 U$$165/A2 U$$14/A1 U$$165/B2 VGND VGND VPWR VPWR U$$150/A sky130_fd_sc_hd__a22o_1
XFILLER_72_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_391_ _407_/CLK _391_/D VGND VGND VPWR VPWR _391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk _380_/CLK VGND VGND VPWR VPWR _397_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_154_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1005 U$$3356/A1 VGND VGND VPWR VPWR U$$4176/B1 sky130_fd_sc_hd__buf_4
XFILLER_193_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1016 U$$477/A1 VGND VGND VPWR VPWR U$$66/A1 sky130_fd_sc_hd__buf_4
XFILLER_5_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1027 U$$3215/A1 VGND VGND VPWR VPWR U$$3213/B1 sky130_fd_sc_hd__buf_6
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1038 U$$3761/A1 VGND VGND VPWR VPWR U$$4309/A1 sky130_fd_sc_hd__buf_6
XFILLER_154_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1049 U$$741/B1 VGND VGND VPWR VPWR U$$878/B1 sky130_fd_sc_hd__buf_4
XFILLER_141_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_74_1 U$$1086/X U$$1219/X U$$1352/X VGND VGND VPWR VPWR dadda_fa_1_75_8/A
+ dadda_fa_1_74_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput240 c[85] VGND VGND VPWR VPWR input240/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_51_0 dadda_fa_3_51_0/A dadda_fa_3_51_0/B dadda_fa_3_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_0/B dadda_fa_4_51_1/CIN sky130_fd_sc_hd__fa_1
Xinput251 c[95] VGND VGND VPWR VPWR input251/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_0_67_0 U$$136/Y U$$273/Y U$$407/X VGND VGND VPWR VPWR dadda_fa_1_68_5/B
+ dadda_fa_1_67_7/B sky130_fd_sc_hd__fa_1
XTAP_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$650 U$$650/A1 U$$652/A2 U$$652/A1 U$$652/B2 VGND VGND VPWR VPWR U$$651/A sky130_fd_sc_hd__a22o_1
XU$$661 U$$661/A U$$684/A VGND VGND VPWR VPWR U$$661/X sky130_fd_sc_hd__xor2_1
XFILLER_17_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$672 U$$807/B1 U$$672/A2 U$$674/A1 U$$553/X VGND VGND VPWR VPWR U$$673/A sky130_fd_sc_hd__a22o_1
XFILLER_17_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$683 U$$683/A U$$683/B VGND VGND VPWR VPWR U$$683/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$694 U$$694/A U$$712/B VGND VGND VPWR VPWR U$$694/X sky130_fd_sc_hd__xor2_1
XFILLER_205_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_11_clk _227_/CLK VGND VGND VPWR VPWR _351_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_96_2 U$$3258/X U$$3391/X U$$3524/X VGND VGND VPWR VPWR dadda_fa_3_97_1/A
+ dadda_fa_3_96_3/A sky130_fd_sc_hd__fa_1
XFILLER_145_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1550 U$$3960/A1 VGND VGND VPWR VPWR U$$4369/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_73_1 dadda_fa_5_73_1/A dadda_fa_5_73_1/B dadda_fa_5_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_74_0/B dadda_fa_7_73_0/A sky130_fd_sc_hd__fa_1
Xrepeater1561 U$$4095/A1 VGND VGND VPWR VPWR U$$4506/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_89_1 U$$3776/X U$$3909/X U$$4042/X VGND VGND VPWR VPWR dadda_fa_3_90_0/CIN
+ dadda_fa_3_89_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater1572 U$$3817/A1 VGND VGND VPWR VPWR U$$3680/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_125_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1583 U$$2582/A1 VGND VGND VPWR VPWR U$$936/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_193_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_66_0 dadda_fa_5_66_0/A dadda_fa_5_66_0/B dadda_fa_5_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_67_0/A dadda_fa_6_66_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1594 input113/X VGND VGND VPWR VPWR U$$4498/A1 sky130_fd_sc_hd__buf_4
XFILLER_154_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_65_8 dadda_fa_1_65_8/A dadda_fa_1_65_8/B dadda_fa_1_65_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_66_3/A dadda_fa_3_65_0/A sky130_fd_sc_hd__fa_2
XFILLER_189_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_58_7 dadda_fa_1_58_7/A dadda_fa_1_58_7/B dadda_fa_1_58_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_59_2/CIN dadda_fa_2_58_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_814 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_5_0 U$$283/X input212/X dadda_fa_6_5_0/CIN VGND VGND VPWR VPWR dadda_fa_7_6_0/B
+ dadda_fa_7_5_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2090 U$$2090/A U$$2092/B VGND VGND VPWR VPWR U$$2090/X sky130_fd_sc_hd__xor2_1
XFILLER_35_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4459_1806 VGND VGND VPWR VPWR U$$4459_1806/HI U$$4459/B sky130_fd_sc_hd__conb_1
XFILLER_50_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_91_1 U$$2317/X U$$2450/X U$$2583/X VGND VGND VPWR VPWR dadda_fa_2_92_4/CIN
+ dadda_fa_2_91_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_84_0 dadda_fa_1_84_0/A U$$1505/X U$$1638/X VGND VGND VPWR VPWR dadda_fa_2_85_2/A
+ dadda_fa_2_84_4/A sky130_fd_sc_hd__fa_1
XFILLER_81_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4409 U$$4409/A U$$4409/B VGND VGND VPWR VPWR U$$4409/X sky130_fd_sc_hd__xor2_1
XTAP_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3708 U$$3708/A U$$3794/B VGND VGND VPWR VPWR U$$3708/X sky130_fd_sc_hd__xor2_1
XFILLER_161_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3719 U$$3719/A1 U$$3739/A2 U$$4269/A1 U$$3739/B2 VGND VGND VPWR VPWR U$$3720/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_374_ _376_/CLK _374_/D VGND VGND VPWR VPWR _374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_83_0 dadda_fa_6_83_0/A dadda_fa_6_83_0/B dadda_fa_6_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_84_0/B dadda_fa_7_83_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_99_0 U$$4461/X input255/X dadda_fa_3_99_0/CIN VGND VGND VPWR VPWR dadda_fa_4_100_0/B
+ dadda_fa_4_99_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$480 U$$480/A U$$484/B VGND VGND VPWR VPWR U$$480/X sky130_fd_sc_hd__xor2_1
XFILLER_211_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$491 U$$763/B1 U$$491/A2 U$$630/A1 U$$491/B2 VGND VGND VPWR VPWR U$$492/A sky130_fd_sc_hd__a22o_1
XFILLER_189_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1380 U$$750/B VGND VGND VPWR VPWR U$$740/B sky130_fd_sc_hd__buf_6
Xrepeater1391 U$$2466/A VGND VGND VPWR VPWR U$$2454/B sky130_fd_sc_hd__buf_8
XFILLER_119_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_70_6 dadda_fa_1_70_6/A dadda_fa_1_70_6/B dadda_fa_1_70_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_2/B dadda_fa_2_70_5/B sky130_fd_sc_hd__fa_1
XFILLER_113_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_63_5 input216/X dadda_fa_1_63_5/B dadda_fa_1_63_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_64_2/A dadda_fa_2_63_5/A sky130_fd_sc_hd__fa_1
XFILLER_41_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_56_4 U$$2779/X U$$2912/X U$$3045/X VGND VGND VPWR VPWR dadda_fa_2_57_1/CIN
+ dadda_fa_2_56_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_49_3 U$$1302/X U$$1435/X U$$1568/X VGND VGND VPWR VPWR dadda_fa_2_50_1/CIN
+ dadda_fa_2_49_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_26_2 dadda_fa_4_26_2/A dadda_fa_4_26_2/B dadda_fa_4_26_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_27_0/CIN dadda_fa_5_26_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_1 dadda_fa_4_19_1/A dadda_fa_4_19_1/B dadda_fa_4_19_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_20_0/B dadda_fa_5_19_1/B sky130_fd_sc_hd__fa_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1085 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4513_1833 VGND VGND VPWR VPWR U$$4513_1833/HI U$$4513/B sky130_fd_sc_hd__conb_1
XFILLER_46_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4206 U$$4478/B1 U$$4210/A2 U$$4343/B1 U$$4210/B2 VGND VGND VPWR VPWR U$$4207/A
+ sky130_fd_sc_hd__a22o_1
XU$$4217 U$$4217/A U$$4247/A VGND VGND VPWR VPWR U$$4217/X sky130_fd_sc_hd__xor2_1
XFILLER_133_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4228 U$$4228/A1 U$$4238/A2 U$$4365/B1 U$$4238/B2 VGND VGND VPWR VPWR U$$4229/A
+ sky130_fd_sc_hd__a22o_1
XU$$4239 U$$4239/A U$$4239/B VGND VGND VPWR VPWR U$$4239/X sky130_fd_sc_hd__xor2_1
XU$$3505 U$$3642/A1 U$$3429/X U$$3644/A1 U$$3430/X VGND VGND VPWR VPWR U$$3506/A sky130_fd_sc_hd__a22o_1
XU$$3516 U$$3516/A U$$3518/B VGND VGND VPWR VPWR U$$3516/X sky130_fd_sc_hd__xor2_1
XU$$3527 U$$4210/B1 U$$3527/A2 U$$3801/B1 U$$3527/B2 VGND VGND VPWR VPWR U$$3528/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3538 U$$3538/A U$$3561/A VGND VGND VPWR VPWR U$$3538/X sky130_fd_sc_hd__xor2_1
XFILLER_45_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3549 U$$3960/A1 U$$3549/A2 U$$3960/B1 U$$3549/B2 VGND VGND VPWR VPWR U$$3550/A
+ sky130_fd_sc_hd__a22o_1
XU$$2804 U$$3352/A1 U$$2810/A2 U$$3078/B1 U$$2810/B2 VGND VGND VPWR VPWR U$$2805/A
+ sky130_fd_sc_hd__a22o_1
XU$$2815 U$$2815/A U$$2817/B VGND VGND VPWR VPWR U$$2815/X sky130_fd_sc_hd__xor2_1
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2826 U$$3511/A1 U$$2874/A2 U$$3648/B1 U$$2874/B2 VGND VGND VPWR VPWR U$$2827/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2837 U$$2837/A U$$2837/B VGND VGND VPWR VPWR U$$2837/X sky130_fd_sc_hd__xor2_1
XANTENNA_120 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2848 U$$2848/A1 U$$2874/A2 U$$4494/A1 U$$2874/B2 VGND VGND VPWR VPWR U$$2849/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _388_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_3_21_1 U$$448/X U$$581/X U$$714/X VGND VGND VPWR VPWR dadda_fa_4_22_0/CIN
+ dadda_fa_4_21_2/A sky130_fd_sc_hd__fa_1
XFILLER_73_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2859 U$$2859/A U$$2859/B VGND VGND VPWR VPWR U$$2859/X sky130_fd_sc_hd__xor2_1
XANTENNA_142 U$$2052/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_153 U$$2828/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_186 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1076 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1038 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_357_ _357_/CLK _357_/D VGND VGND VPWR VPWR _357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_288_ _417_/CLK _288_/D VGND VGND VPWR VPWR _288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_80_5 dadda_fa_2_80_5/A dadda_fa_2_80_5/B dadda_fa_2_80_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_81_2/A dadda_fa_4_80_0/A sky130_fd_sc_hd__fa_2
XFILLER_68_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_73_4 dadda_fa_2_73_4/A dadda_fa_2_73_4/B dadda_fa_2_73_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_1/CIN dadda_fa_3_73_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_66_3 dadda_fa_2_66_3/A dadda_fa_2_66_3/B dadda_fa_2_66_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/B dadda_fa_3_66_3/B sky130_fd_sc_hd__fa_2
XFILLER_68_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_59_2 dadda_fa_2_59_2/A dadda_fa_2_59_2/B dadda_fa_2_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/A dadda_fa_3_59_3/A sky130_fd_sc_hd__fa_1
XFILLER_83_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 a[12] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_1083 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_36_1 dadda_fa_5_36_1/A dadda_fa_5_36_1/B dadda_fa_5_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_37_0/B dadda_fa_7_36_0/A sky130_fd_sc_hd__fa_1
XFILLER_65_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_29_0 dadda_fa_5_29_0/A dadda_fa_5_29_0/B dadda_fa_5_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_30_0/A dadda_fa_6_29_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_36_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_110_1 dadda_fa_5_110_1/A dadda_fa_5_110_1/B dadda_fa_5_110_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_111_0/B dadda_fa_7_110_0/A sky130_fd_sc_hd__fa_1
XFILLER_192_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$2 _298_/Q _170_/Q VGND VGND VPWR VPWR final_adder.U$$253/A2 final_adder.U$$252/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_5_103_0 dadda_fa_5_103_0/A dadda_fa_5_103_0/B dadda_fa_5_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_104_0/A dadda_fa_6_103_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_106_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput330 output330/A VGND VGND VPWR VPWR o[50] sky130_fd_sc_hd__buf_2
XFILLER_10_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput341 output341/A VGND VGND VPWR VPWR o[60] sky130_fd_sc_hd__buf_2
XFILLER_156_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput352 output352/A VGND VGND VPWR VPWR o[70] sky130_fd_sc_hd__buf_2
XFILLER_0_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput363 output363/A VGND VGND VPWR VPWR o[80] sky130_fd_sc_hd__buf_2
Xoutput374 output374/A VGND VGND VPWR VPWR o[90] sky130_fd_sc_hd__buf_2
XFILLER_114_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_671 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_61_2 U$$2789/X U$$2922/X U$$3055/X VGND VGND VPWR VPWR dadda_fa_2_62_1/A
+ dadda_fa_2_61_4/A sky130_fd_sc_hd__fa_1
XFILLER_142_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_54_1 U$$1179/X U$$1312/X U$$1445/X VGND VGND VPWR VPWR dadda_fa_2_55_0/CIN
+ dadda_fa_2_54_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_31_0 dadda_fa_4_31_0/A dadda_fa_4_31_0/B dadda_fa_4_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/A dadda_fa_5_31_1/A sky130_fd_sc_hd__fa_1
XFILLER_90_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_47_0 U$$101/X U$$234/X U$$367/X VGND VGND VPWR VPWR dadda_fa_2_48_1/B
+ dadda_fa_2_47_4/A sky130_fd_sc_hd__fa_1
XFILLER_83_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_211_ _211_/CLK _211_/D VGND VGND VPWR VPWR _211_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_208_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_83_3 dadda_fa_3_83_3/A dadda_fa_3_83_3/B dadda_fa_3_83_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_84_1/B dadda_fa_4_83_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_76_2 dadda_fa_3_76_2/A dadda_fa_3_76_2/B dadda_fa_3_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_1/A dadda_fa_4_76_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_3_69_1 dadda_fa_3_69_1/A dadda_fa_3_69_1/B dadda_fa_3_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_0/CIN dadda_fa_4_69_2/A sky130_fd_sc_hd__fa_1
XFILLER_78_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_46_0 dadda_fa_6_46_0/A dadda_fa_6_46_0/B dadda_fa_6_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_47_0/B dadda_fa_7_46_0/CIN sky130_fd_sc_hd__fa_1
XU$$4003 U$$4275/B1 U$$4035/A2 U$$4277/B1 U$$4035/B2 VGND VGND VPWR VPWR U$$4004/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4014 U$$4014/A U$$4080/B VGND VGND VPWR VPWR U$$4014/X sky130_fd_sc_hd__xor2_1
XU$$4025 U$$4162/A1 U$$4043/A2 U$$4162/B1 U$$4043/B2 VGND VGND VPWR VPWR U$$4026/A
+ sky130_fd_sc_hd__a22o_1
XU$$4036 U$$4036/A U$$4036/B VGND VGND VPWR VPWR U$$4036/X sky130_fd_sc_hd__xor2_1
XFILLER_59_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3302 U$$3713/A1 U$$3394/A2 U$$3578/A1 U$$3394/B2 VGND VGND VPWR VPWR U$$3303/A
+ sky130_fd_sc_hd__a22o_1
XU$$3422_1748 VGND VGND VPWR VPWR U$$3422_1748/HI U$$3422/B1 sky130_fd_sc_hd__conb_1
XFILLER_93_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4047 input91/X U$$4107/A2 input92/X U$$4107/B2 VGND VGND VPWR VPWR U$$4048/A sky130_fd_sc_hd__a22o_1
XFILLER_111_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4058 U$$4058/A U$$4078/B VGND VGND VPWR VPWR U$$4058/X sky130_fd_sc_hd__xor2_1
XU$$3313 U$$3313/A U$$3349/B VGND VGND VPWR VPWR U$$3313/X sky130_fd_sc_hd__xor2_1
XFILLER_47_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4069 input103/X U$$4079/A2 input104/X U$$4079/B2 VGND VGND VPWR VPWR U$$4070/A
+ sky130_fd_sc_hd__a22o_1
XU$$3324 U$$4009/A1 U$$3348/A2 U$$860/A1 U$$3346/B2 VGND VGND VPWR VPWR U$$3325/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3335 U$$3335/A U$$3375/B VGND VGND VPWR VPWR U$$3335/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_1211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2601 U$$2601/A U$$2601/B VGND VGND VPWR VPWR U$$2601/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3346 U$$741/B1 U$$3348/A2 U$$3485/A1 U$$3346/B2 VGND VGND VPWR VPWR U$$3347/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2612 U$$2612/A U$$2624/B VGND VGND VPWR VPWR U$$2612/X sky130_fd_sc_hd__xor2_1
XFILLER_206_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_105_2 dadda_fa_4_105_2/A dadda_fa_4_105_2/B dadda_fa_4_105_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_106_0/CIN dadda_fa_5_105_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_20_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3357 U$$3357/A U$$3389/B VGND VGND VPWR VPWR U$$3357/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3368 U$$3642/A1 U$$3374/A2 U$$3368/B1 U$$3374/B2 VGND VGND VPWR VPWR U$$3369/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2623 U$$2623/A1 U$$2625/A2 U$$2625/A1 U$$2625/B2 VGND VGND VPWR VPWR U$$2624/A
+ sky130_fd_sc_hd__a22o_1
XU$$2634 U$$2634/A U$$2650/B VGND VGND VPWR VPWR U$$2634/X sky130_fd_sc_hd__xor2_1
XFILLER_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3379 U$$3379/A U$$3425/A VGND VGND VPWR VPWR U$$3379/X sky130_fd_sc_hd__xor2_1
XU$$2645 U$$4013/B1 U$$2727/A2 U$$4015/B1 U$$2727/B2 VGND VGND VPWR VPWR U$$2646/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1900 U$$1900/A U$$1914/B VGND VGND VPWR VPWR U$$1900/X sky130_fd_sc_hd__xor2_1
XU$$1911 U$$4514/A1 U$$1785/X U$$4516/A1 U$$1786/X VGND VGND VPWR VPWR U$$1912/A sky130_fd_sc_hd__a22o_1
XU$$2656 U$$2656/A U$$2658/B VGND VGND VPWR VPWR U$$2656/X sky130_fd_sc_hd__xor2_1
XFILLER_206_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2667 U$$3352/A1 U$$2607/X U$$3078/B1 U$$2608/X VGND VGND VPWR VPWR U$$2668/A sky130_fd_sc_hd__a22o_1
XU$$1922 U$$1920/Y input21/X input20/X U$$1921/X U$$1918/Y VGND VGND VPWR VPWR U$$1922/X
+ sky130_fd_sc_hd__a32o_2
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1933 U$$1933/A U$$1971/B VGND VGND VPWR VPWR U$$1933/X sky130_fd_sc_hd__xor2_1
XU$$2678 U$$2678/A U$$2680/B VGND VGND VPWR VPWR U$$2678/X sky130_fd_sc_hd__xor2_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2689 U$$4468/B1 U$$2737/A2 U$$3648/B1 U$$2737/B2 VGND VGND VPWR VPWR U$$2690/A
+ sky130_fd_sc_hd__a22o_1
XU$$1944 U$$2492/A1 U$$1960/A2 U$$3453/A1 U$$1960/B2 VGND VGND VPWR VPWR U$$1945/A
+ sky130_fd_sc_hd__a22o_1
XU$$1955 U$$1955/A U$$1993/B VGND VGND VPWR VPWR U$$1955/X sky130_fd_sc_hd__xor2_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1966 U$$3747/A1 U$$1970/A2 U$$50/A1 U$$1970/B2 VGND VGND VPWR VPWR U$$1967/A sky130_fd_sc_hd__a22o_1
XFILLER_199_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1977 U$$1977/A U$$2017/B VGND VGND VPWR VPWR U$$1977/X sky130_fd_sc_hd__xor2_1
XFILLER_15_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1988 U$$616/B1 U$$1990/A2 U$$2810/B1 U$$1990/B2 VGND VGND VPWR VPWR U$$1989/A
+ sky130_fd_sc_hd__a22o_1
X_409_ _411_/CLK _409_/D VGND VGND VPWR VPWR _409_/Q sky130_fd_sc_hd__dfxtp_1
XU$$1999 U$$1999/A U$$2043/B VGND VGND VPWR VPWR U$$1999/X sky130_fd_sc_hd__xor2_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_119_0 dadda_fa_7_119_0/A dadda_fa_7_119_0/B dadda_fa_7_119_0/CIN VGND
+ VGND VPWR VPWR _416_/D _287_/D sky130_fd_sc_hd__fa_1
XFILLER_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_71_1 dadda_fa_2_71_1/A dadda_fa_2_71_1/B dadda_fa_2_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_0/CIN dadda_fa_3_71_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_64_0 dadda_fa_2_64_0/A dadda_fa_2_64_0/B dadda_fa_2_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_0/B dadda_fa_3_64_2/B sky130_fd_sc_hd__fa_1
XFILLER_97_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater800 U$$2334/X VGND VGND VPWR VPWR U$$2403/B2 sky130_fd_sc_hd__clkbuf_8
Xfinal_adder.U$$607 final_adder.U$$606/B final_adder.U$$491/X final_adder.U$$483/X
+ VGND VGND VPWR VPWR final_adder.U$$607/X sky130_fd_sc_hd__a21o_1
XFILLER_69_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater811 U$$2316/B2 VGND VGND VPWR VPWR U$$2326/B2 sky130_fd_sc_hd__buf_4
XFILLER_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater822 U$$2060/X VGND VGND VPWR VPWR U$$2177/B2 sky130_fd_sc_hd__buf_6
XFILLER_111_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$629 final_adder.U$$628/B final_adder.U$$525/X final_adder.U$$509/X
+ VGND VGND VPWR VPWR final_adder.U$$629/X sky130_fd_sc_hd__a21o_1
XFILLER_38_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater833 U$$1903/B2 VGND VGND VPWR VPWR U$$1879/B2 sky130_fd_sc_hd__buf_4
Xrepeater844 U$$1770/B2 VGND VGND VPWR VPWR U$$1764/B2 sky130_fd_sc_hd__buf_6
XFILLER_110_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater855 U$$231/B2 VGND VGND VPWR VPWR U$$217/B2 sky130_fd_sc_hd__buf_6
Xrepeater866 U$$1470/B2 VGND VGND VPWR VPWR U$$1422/B2 sky130_fd_sc_hd__buf_4
XFILLER_42_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater877 U$$1337/B2 VGND VGND VPWR VPWR U$$1291/B2 sky130_fd_sc_hd__buf_4
Xrepeater888 U$$42/B2 VGND VGND VPWR VPWR U$$8/B2 sky130_fd_sc_hd__buf_4
Xrepeater899 U$$4494/B2 VGND VGND VPWR VPWR U$$4486/B2 sky130_fd_sc_hd__clkbuf_4
XU$$40 U$$40/A1 U$$42/A2 U$$42/A1 U$$42/B2 VGND VGND VPWR VPWR U$$41/A sky130_fd_sc_hd__a22o_1
XFILLER_71_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$51 U$$51/A U$$51/B VGND VGND VPWR VPWR U$$51/X sky130_fd_sc_hd__xor2_1
XU$$62 U$$62/A1 U$$94/A2 U$$62/B1 U$$94/B2 VGND VGND VPWR VPWR U$$63/A sky130_fd_sc_hd__a22o_1
XFILLER_53_923 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$73 U$$73/A U$$81/B VGND VGND VPWR VPWR U$$73/X sky130_fd_sc_hd__xor2_1
XU$$84 U$$84/A1 U$$98/A2 U$$84/B1 U$$98/B2 VGND VGND VPWR VPWR U$$85/A sky130_fd_sc_hd__a22o_1
XU$$3880 input74/X U$$3970/A2 U$$3880/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3881/A
+ sky130_fd_sc_hd__a22o_1
XU$$95 U$$95/A U$$99/B VGND VGND VPWR VPWR U$$95/X sky130_fd_sc_hd__xor2_1
XFILLER_52_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3891 U$$3891/A U$$3909/B VGND VGND VPWR VPWR U$$3891/X sky130_fd_sc_hd__xor2_1
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1055 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_20 _336_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_31 _339_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_42 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _342_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_75 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_86 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_97 _346_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_4_93_2 dadda_fa_4_93_2/A dadda_fa_4_93_2/B dadda_fa_4_93_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_94_0/CIN dadda_fa_5_93_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_86_1 dadda_fa_4_86_1/A dadda_fa_4_86_1/B dadda_fa_4_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/B dadda_fa_5_86_1/B sky130_fd_sc_hd__fa_1
XFILLER_161_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_63_0 dadda_fa_7_63_0/A dadda_fa_7_63_0/B dadda_fa_7_63_0/CIN VGND VGND
+ VPWR VPWR _360_/D _231_/D sky130_fd_sc_hd__fa_1
XFILLER_133_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_79_0 dadda_fa_4_79_0/A dadda_fa_4_79_0/B dadda_fa_4_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/A dadda_fa_5_79_1/A sky130_fd_sc_hd__fa_1
XFILLER_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1075 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1207 U$$1207/A U$$1209/B VGND VGND VPWR VPWR U$$1207/X sky130_fd_sc_hd__xor2_1
XFILLER_55_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1218 U$$944/A1 U$$1230/A2 U$$944/B1 U$$1230/B2 VGND VGND VPWR VPWR U$$1219/A sky130_fd_sc_hd__a22o_1
XFILLER_189_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1229 U$$1229/A U$$1232/A VGND VGND VPWR VPWR U$$1229/X sky130_fd_sc_hd__xor2_1
XFILLER_203_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1001 final_adder.U$$230/A final_adder.U$$731/X final_adder.U$$231/A2
+ VGND VGND VPWR VPWR final_adder.U$$1049/B sky130_fd_sc_hd__a21o_1
XFILLER_200_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1023 final_adder.U$$252/A final_adder.U$$255/X final_adder.U$$253/A2
+ VGND VGND VPWR VPWR final_adder.U$$1027/B sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$1034 final_adder.U$$244/A final_adder.U$$625/X VGND VGND VPWR VPWR
+ output268/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1045 final_adder.U$$234/B final_adder.U$$1045/B VGND VGND VPWR VPWR
+ output298/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1056 final_adder.U$$222/A final_adder.U$$723/X VGND VGND VPWR VPWR
+ output310/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1067 final_adder.U$$212/B final_adder.U$$983/X VGND VGND VPWR VPWR
+ output322/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1078 final_adder.U$$200/A final_adder.U$$813/X VGND VGND VPWR VPWR
+ output334/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1089 final_adder.U$$190/B final_adder.U$$961/X VGND VGND VPWR VPWR
+ output346/A sky130_fd_sc_hd__xor2_1
XFILLER_125_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_81_0 dadda_fa_3_81_0/A dadda_fa_3_81_0/B dadda_fa_3_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_0/B dadda_fa_4_81_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_125_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_396 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3110 U$$3245/B1 U$$3018/X U$$3112/A1 U$$3019/X VGND VGND VPWR VPWR U$$3111/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_110_0 input141/X dadda_fa_4_110_0/B dadda_fa_4_110_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_5_111_0/A dadda_fa_5_110_1/A sky130_fd_sc_hd__fa_1
XU$$3121 U$$3121/A U$$3133/B VGND VGND VPWR VPWR U$$3121/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_43_5 dadda_fa_2_43_5/A dadda_fa_2_43_5/B dadda_fa_2_43_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_44_2/A dadda_fa_4_43_0/A sky130_fd_sc_hd__fa_2
XFILLER_4_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3132 U$$3680/A1 U$$3132/A2 U$$118/B1 U$$3132/B2 VGND VGND VPWR VPWR U$$3133/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3143 U$$3143/A U$$3150/A VGND VGND VPWR VPWR U$$3143/X sky130_fd_sc_hd__xor2_1
XFILLER_207_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3154 U$$3288/A U$$3154/B VGND VGND VPWR VPWR U$$3154/X sky130_fd_sc_hd__and2_1
XU$$2420 U$$2420/A U$$2465/A VGND VGND VPWR VPWR U$$2420/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_36_4 U$$2340/X U$$2473/X U$$2525/B VGND VGND VPWR VPWR dadda_fa_3_37_1/CIN
+ dadda_fa_3_36_3/CIN sky130_fd_sc_hd__fa_1
XU$$3165 U$$3300/B1 U$$3187/A2 input109/X U$$3187/B2 VGND VGND VPWR VPWR U$$3166/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2431 U$$3116/A1 U$$2333/X U$$3116/B1 U$$2334/X VGND VGND VPWR VPWR U$$2432/A sky130_fd_sc_hd__a22o_1
XFILLER_185_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3176 U$$3176/A U$$3264/B VGND VGND VPWR VPWR U$$3176/X sky130_fd_sc_hd__xor2_1
XU$$2442 U$$2442/A U$$2442/B VGND VGND VPWR VPWR U$$2442/X sky130_fd_sc_hd__xor2_1
XU$$3187 U$$4144/B1 U$$3187/A2 U$$4422/A1 U$$3187/B2 VGND VGND VPWR VPWR U$$3188/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2453 U$$3960/A1 U$$2459/A2 U$$3960/B1 U$$2459/B2 VGND VGND VPWR VPWR U$$2454/A
+ sky130_fd_sc_hd__a22o_1
XU$$3198 U$$3198/A U$$3242/B VGND VGND VPWR VPWR U$$3198/X sky130_fd_sc_hd__xor2_1
XU$$2464 U$$2464/A U$$2465/A VGND VGND VPWR VPWR U$$2464/X sky130_fd_sc_hd__xor2_1
XFILLER_50_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1730 U$$2415/A1 U$$1736/A2 U$$2691/A1 U$$1736/B2 VGND VGND VPWR VPWR U$$1731/A
+ sky130_fd_sc_hd__a22o_1
XU$$2475 U$$2475/A U$$2525/B VGND VGND VPWR VPWR U$$2475/X sky130_fd_sc_hd__xor2_1
XU$$2486 U$$2623/A1 U$$2490/A2 U$$2625/A1 U$$2490/B2 VGND VGND VPWR VPWR U$$2487/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1741 U$$1741/A U$$1780/A VGND VGND VPWR VPWR U$$1741/X sky130_fd_sc_hd__xor2_1
XFILLER_62_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1752 U$$517/B1 U$$1764/A2 U$$384/A1 U$$1764/B2 VGND VGND VPWR VPWR U$$1753/A sky130_fd_sc_hd__a22o_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2497 U$$2497/A U$$2543/B VGND VGND VPWR VPWR U$$2497/X sky130_fd_sc_hd__xor2_1
XU$$1763 U$$1763/A U$$1765/B VGND VGND VPWR VPWR U$$1763/X sky130_fd_sc_hd__xor2_1
XU$$1774 U$$4514/A1 U$$1648/X U$$4516/A1 U$$1649/X VGND VGND VPWR VPWR U$$1775/A sky130_fd_sc_hd__a22o_1
XU$$1785 U$$1783/Y input19/X input18/X U$$1784/X U$$1781/Y VGND VGND VPWR VPWR U$$1785/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_21_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1796 U$$1796/A U$$1832/B VGND VGND VPWR VPWR U$$1796/X sky130_fd_sc_hd__xor2_1
XFILLER_175_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_96_0 dadda_fa_5_96_0/A dadda_fa_5_96_0/B dadda_fa_5_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_97_0/A dadda_fa_6_96_0/CIN sky130_fd_sc_hd__fa_1
Xinput40 a[45] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput51 a[55] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput62 a[7] VGND VGND VPWR VPWR U$$548/A sky130_fd_sc_hd__buf_6
XFILLER_162_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput73 b[17] VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__buf_8
Xinput84 b[27] VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__buf_8
Xinput95 b[37] VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__buf_8
XFILLER_190_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$404 final_adder.U$$408/B final_adder.U$$404/B VGND VGND VPWR VPWR
+ final_adder.U$$528/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$415 final_adder.U$$414/B final_adder.U$$293/X final_adder.U$$289/X
+ VGND VGND VPWR VPWR final_adder.U$$415/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$426 final_adder.U$$430/B final_adder.U$$426/B VGND VGND VPWR VPWR
+ final_adder.U$$550/B sky130_fd_sc_hd__and2_1
Xrepeater630 U$$1237/X VGND VGND VPWR VPWR U$$1353/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$437 final_adder.U$$436/B final_adder.U$$315/X final_adder.U$$311/X
+ VGND VGND VPWR VPWR final_adder.U$$437/X sky130_fd_sc_hd__a21o_1
XTAP_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater641 U$$997/B2 VGND VGND VPWR VPWR U$$999/B2 sky130_fd_sc_hd__buf_4
XFILLER_85_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$448 final_adder.U$$452/B final_adder.U$$448/B VGND VGND VPWR VPWR
+ final_adder.U$$572/B sky130_fd_sc_hd__and2_1
XTAP_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater652 U$$950/B2 VGND VGND VPWR VPWR U$$918/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$459 final_adder.U$$458/B final_adder.U$$337/X final_adder.U$$333/X
+ VGND VGND VPWR VPWR final_adder.U$$459/X sky130_fd_sc_hd__a21o_1
Xrepeater663 U$$668/B2 VGND VGND VPWR VPWR U$$624/B2 sky130_fd_sc_hd__buf_4
Xrepeater674 U$$4361/B2 VGND VGND VPWR VPWR U$$4349/B2 sky130_fd_sc_hd__clkbuf_4
XU$$309 U$$309/A U$$317/B VGND VGND VPWR VPWR U$$309/X sky130_fd_sc_hd__xor2_1
Xrepeater685 U$$416/X VGND VGND VPWR VPWR U$$537/B2 sky130_fd_sc_hd__buf_6
Xrepeater696 U$$4079/B2 VGND VGND VPWR VPWR U$$4077/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1209 U$$683/B VGND VGND VPWR VPWR U$$684/A sky130_fd_sc_hd__buf_8
XFILLER_181_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_105_1 U$$4074/X U$$4207/X U$$4340/X VGND VGND VPWR VPWR dadda_fa_4_106_0/CIN
+ dadda_fa_4_105_2/A sky130_fd_sc_hd__fa_1
XFILLER_106_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_126_0 U$$4515/X input158/X dadda_fa_6_126_0/CIN VGND VGND VPWR VPWR dadda_fa_7_127_0/B
+ dadda_fa_7_126_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_69_4 U$$2007/X U$$2140/X U$$2273/X VGND VGND VPWR VPWR dadda_fa_1_70_7/B
+ dadda_fa_2_69_0/A sky130_fd_sc_hd__fa_1
XTAP_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_46_3 dadda_fa_3_46_3/A dadda_fa_3_46_3/B dadda_fa_3_46_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_47_1/B dadda_fa_4_46_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$971 final_adder.U$$200/A final_adder.U$$813/X final_adder.U$$971/B1
+ VGND VGND VPWR VPWR final_adder.U$$971/X sky130_fd_sc_hd__a21o_1
XU$$810 U$$810/A U$$821/A VGND VGND VPWR VPWR U$$810/X sky130_fd_sc_hd__xor2_1
XFILLER_63_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_39_2 dadda_fa_3_39_2/A dadda_fa_3_39_2/B dadda_fa_3_39_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_1/A dadda_fa_4_39_2/B sky130_fd_sc_hd__fa_1
XU$$821 U$$821/A VGND VGND VPWR VPWR U$$821/Y sky130_fd_sc_hd__inv_1
XTAP_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$993 final_adder.U$$222/A final_adder.U$$723/X final_adder.U$$993/B1
+ VGND VGND VPWR VPWR final_adder.U$$993/X sky130_fd_sc_hd__a21o_1
XU$$832 U$$832/A1 U$$918/A2 U$$969/B1 U$$918/B2 VGND VGND VPWR VPWR U$$833/A sky130_fd_sc_hd__a22o_1
XFILLER_44_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_4_122_0_1875 VGND VGND VPWR VPWR dadda_ha_4_122_0/A dadda_ha_4_122_0_1875/LO
+ sky130_fd_sc_hd__conb_1
XU$$843 U$$843/A U$$847/B VGND VGND VPWR VPWR U$$843/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$854 U$$854/A1 U$$882/A2 U$$854/B1 U$$882/B2 VGND VGND VPWR VPWR U$$855/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$865 U$$865/A U$$883/B VGND VGND VPWR VPWR U$$865/X sky130_fd_sc_hd__xor2_1
XU$$1004 U$$1004/A U$$996/B VGND VGND VPWR VPWR U$$1004/X sky130_fd_sc_hd__xor2_1
XU$$1015 U$$330/A1 U$$997/A2 U$$56/B1 U$$997/B2 VGND VGND VPWR VPWR U$$1016/A sky130_fd_sc_hd__a22o_1
XU$$876 U$$54/A1 U$$882/A2 U$$56/A1 U$$882/B2 VGND VGND VPWR VPWR U$$877/A sky130_fd_sc_hd__a22o_1
XU$$1026 U$$1026/A U$$994/B VGND VGND VPWR VPWR U$$1026/X sky130_fd_sc_hd__xor2_1
XFILLER_73_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$887 U$$887/A U$$929/B VGND VGND VPWR VPWR U$$887/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$898 U$$76/A1 U$$950/A2 U$$78/A1 U$$950/B2 VGND VGND VPWR VPWR U$$899/A sky130_fd_sc_hd__a22o_1
XFILLER_91_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1037 U$$1448/A1 U$$979/A2 U$$902/A1 U$$979/B2 VGND VGND VPWR VPWR U$$1038/A sky130_fd_sc_hd__a22o_1
XU$$1048 U$$1048/A U$$968/B VGND VGND VPWR VPWR U$$1048/X sky130_fd_sc_hd__xor2_1
XFILLER_16_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_414 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1059 U$$98/B1 U$$1083/A2 U$$924/A1 U$$1083/B2 VGND VGND VPWR VPWR U$$1060/A sky130_fd_sc_hd__a22o_1
XFILLER_31_469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_41_2 U$$2350/X U$$2483/X U$$2616/X VGND VGND VPWR VPWR dadda_fa_3_42_1/A
+ dadda_fa_3_41_3/A sky130_fd_sc_hd__fa_1
XFILLER_148_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_34_1 U$$740/X U$$873/X U$$1006/X VGND VGND VPWR VPWR dadda_fa_3_35_0/CIN
+ dadda_fa_3_34_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_207_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_11_0 U$$694/X input151/X dadda_fa_5_11_0/CIN VGND VGND VPWR VPWR dadda_fa_6_12_0/A
+ dadda_fa_6_11_0/CIN sky130_fd_sc_hd__fa_1
XU$$2250 U$$741/B1 U$$2252/A2 U$$3483/B1 U$$2252/B2 VGND VGND VPWR VPWR U$$2251/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_27_0 U$$61/X U$$194/X U$$327/X VGND VGND VPWR VPWR dadda_fa_3_28_2/A dadda_fa_3_27_3/B
+ sky130_fd_sc_hd__fa_1
XU$$2261 U$$2261/A U$$2309/B VGND VGND VPWR VPWR U$$2261/X sky130_fd_sc_hd__xor2_1
XFILLER_22_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2272 U$$2957/A1 U$$2272/A2 U$$2409/B1 U$$2272/B2 VGND VGND VPWR VPWR U$$2273/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2283 U$$2283/A U$$2303/B VGND VGND VPWR VPWR U$$2283/X sky130_fd_sc_hd__xor2_1
XU$$2294 U$$3116/A1 U$$2316/A2 U$$3116/B1 U$$2316/B2 VGND VGND VPWR VPWR U$$2295/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1560 U$$1560/A U$$1592/B VGND VGND VPWR VPWR U$$1560/X sky130_fd_sc_hd__xor2_1
XU$$1571 U$$3215/A1 U$$1575/A2 U$$1984/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1572/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1582 U$$1582/A U$$1620/B VGND VGND VPWR VPWR U$$1582/X sky130_fd_sc_hd__xor2_1
XU$$1593 U$$86/A1 U$$1607/A2 U$$88/A1 U$$1607/B2 VGND VGND VPWR VPWR U$$1594/A sky130_fd_sc_hd__a22o_1
XFILLER_163_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_86_4 U$$3105/X U$$3238/X U$$3371/X VGND VGND VPWR VPWR dadda_fa_2_87_4/A
+ dadda_fa_2_86_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_104_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_79_3 U$$2293/X U$$2426/X U$$2559/X VGND VGND VPWR VPWR dadda_fa_2_80_1/B
+ dadda_fa_2_79_4/B sky130_fd_sc_hd__fa_1
XFILLER_58_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_56_2 dadda_fa_4_56_2/A dadda_fa_4_56_2/B dadda_fa_4_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_57_0/CIN dadda_fa_5_56_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$201 final_adder.U$$200/B final_adder.U$$971/B1 final_adder.U$$201/B1
+ VGND VGND VPWR VPWR final_adder.U$$201/X sky130_fd_sc_hd__a21o_1
XFILLER_134_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$212 final_adder.U$$212/A final_adder.U$$212/B VGND VGND VPWR VPWR
+ final_adder.U$$340/B sky130_fd_sc_hd__and2_1
XTAP_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$223 final_adder.U$$222/B final_adder.U$$993/B1 final_adder.U$$223/B1
+ VGND VGND VPWR VPWR final_adder.U$$223/X sky130_fd_sc_hd__a21o_1
XTAP_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_49_1 dadda_fa_4_49_1/A dadda_fa_4_49_1/B dadda_fa_4_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/B dadda_fa_5_49_1/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$234 final_adder.U$$234/A final_adder.U$$234/B VGND VGND VPWR VPWR
+ final_adder.U$$362/B sky130_fd_sc_hd__and2_1
XTAP_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$245 final_adder.U$$244/B final_adder.U$$245/A2 final_adder.U$$245/B1
+ VGND VGND VPWR VPWR final_adder.U$$245/X sky130_fd_sc_hd__a21o_1
XTAP_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater460 U$$3966/A2 VGND VGND VPWR VPWR U$$3926/A2 sky130_fd_sc_hd__buf_6
XTAP_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_26_0 dadda_fa_7_26_0/A dadda_fa_7_26_0/B dadda_fa_7_26_0/CIN VGND VGND
+ VPWR VPWR _323_/D _194_/D sky130_fd_sc_hd__fa_2
XFILLER_79_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$267 final_adder.U$$266/B final_adder.U$$141/X final_adder.U$$139/X
+ VGND VGND VPWR VPWR final_adder.U$$267/X sky130_fd_sc_hd__a21o_1
XTAP_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater471 U$$3612/A2 VGND VGND VPWR VPWR U$$3606/A2 sky130_fd_sc_hd__buf_6
XU$$106 U$$654/A1 U$$122/A2 U$$654/B1 U$$122/B2 VGND VGND VPWR VPWR U$$107/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$278 final_adder.U$$280/B final_adder.U$$278/B VGND VGND VPWR VPWR
+ final_adder.U$$404/B sky130_fd_sc_hd__and2_1
XU$$117 U$$117/A U$$127/B VGND VGND VPWR VPWR U$$117/X sky130_fd_sc_hd__xor2_1
XTAP_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater482 U$$3489/A2 VGND VGND VPWR VPWR U$$3527/A2 sky130_fd_sc_hd__buf_6
XFILLER_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$289 final_adder.U$$288/B final_adder.U$$163/X final_adder.U$$161/X
+ VGND VGND VPWR VPWR final_adder.U$$289/X sky130_fd_sc_hd__a21o_1
XU$$128 U$$950/A1 U$$134/A2 U$$676/B1 U$$134/B2 VGND VGND VPWR VPWR U$$129/A sky130_fd_sc_hd__a22o_1
Xrepeater493 U$$3378/A2 VGND VGND VPWR VPWR U$$3388/A2 sky130_fd_sc_hd__buf_6
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$139 U$$272/B VGND VGND VPWR VPWR U$$139/Y sky130_fd_sc_hd__inv_1
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_390_ _390_/CLK _390_/D VGND VGND VPWR VPWR _390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4401_1777 VGND VGND VPWR VPWR U$$4401_1777/HI U$$4401/B sky130_fd_sc_hd__conb_1
XFILLER_175_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1006 input88/X VGND VGND VPWR VPWR U$$3356/A1 sky130_fd_sc_hd__buf_6
XFILLER_181_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1017 U$$1984/A1 VGND VGND VPWR VPWR U$$477/A1 sky130_fd_sc_hd__buf_4
Xrepeater1028 input85/X VGND VGND VPWR VPWR U$$3215/A1 sky130_fd_sc_hd__buf_4
XFILLER_135_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1039 input84/X VGND VGND VPWR VPWR U$$3761/A1 sky130_fd_sc_hd__buf_6
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput230 c[76] VGND VGND VPWR VPWR input230/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_51_1 dadda_fa_3_51_1/A dadda_fa_3_51_1/B dadda_fa_3_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_0/CIN dadda_fa_4_51_2/A sky130_fd_sc_hd__fa_1
Xinput241 c[86] VGND VGND VPWR VPWR input241/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_67_1 U$$540/X U$$673/X U$$806/X VGND VGND VPWR VPWR dadda_fa_1_68_5/CIN
+ dadda_fa_1_67_7/CIN sky130_fd_sc_hd__fa_1
Xinput252 c[96] VGND VGND VPWR VPWR input252/X sky130_fd_sc_hd__clkbuf_4
XTAP_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_44_0 dadda_fa_3_44_0/A dadda_fa_3_44_0/B dadda_fa_3_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_0/B dadda_fa_4_44_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$790 final_adder.U$$790/A final_adder.U$$790/B VGND VGND VPWR VPWR
+ final_adder.U$$790/X sky130_fd_sc_hd__and2_1
XFILLER_29_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$640 U$$640/A1 U$$652/A2 U$$916/A1 U$$652/B2 VGND VGND VPWR VPWR U$$641/A sky130_fd_sc_hd__a22o_1
XFILLER_112_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$651 U$$651/A U$$651/B VGND VGND VPWR VPWR U$$651/X sky130_fd_sc_hd__xor2_1
XU$$662 U$$799/A1 U$$672/A2 U$$938/A1 U$$668/B2 VGND VGND VPWR VPWR U$$663/A sky130_fd_sc_hd__a22o_1
XFILLER_210_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$673 U$$673/A U$$673/B VGND VGND VPWR VPWR U$$673/X sky130_fd_sc_hd__xor2_1
XFILLER_205_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$684 U$$684/A VGND VGND VPWR VPWR U$$684/Y sky130_fd_sc_hd__inv_1
XU$$695 U$$832/A1 U$$783/A2 U$$969/B1 U$$783/B2 VGND VGND VPWR VPWR U$$696/A sky130_fd_sc_hd__a22o_1
XFILLER_17_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_974 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_101_0 dadda_fa_7_101_0/A dadda_fa_7_101_0/B dadda_fa_7_101_0/CIN VGND
+ VGND VPWR VPWR _398_/D _269_/D sky130_fd_sc_hd__fa_1
XFILLER_172_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_96_3 U$$3657/X U$$3790/X U$$3923/X VGND VGND VPWR VPWR dadda_fa_3_97_1/B
+ dadda_fa_3_96_3/B sky130_fd_sc_hd__fa_1
XFILLER_172_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1540 U$$4236/A1 VGND VGND VPWR VPWR U$$811/A1 sky130_fd_sc_hd__buf_4
Xrepeater1551 U$$4508/A1 VGND VGND VPWR VPWR U$$807/B1 sky130_fd_sc_hd__buf_4
XFILLER_67_1143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1562 input117/X VGND VGND VPWR VPWR U$$4095/A1 sky130_fd_sc_hd__buf_4
XFILLER_141_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_89_2 U$$4175/X U$$4308/X U$$4441/X VGND VGND VPWR VPWR dadda_fa_3_90_1/A
+ dadda_fa_3_89_3/A sky130_fd_sc_hd__fa_1
XFILLER_141_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1573 U$$4502/A1 VGND VGND VPWR VPWR U$$527/B1 sky130_fd_sc_hd__buf_6
XFILLER_125_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1584 U$$4500/A1 VGND VGND VPWR VPWR U$$2582/A1 sky130_fd_sc_hd__buf_4
XFILLER_119_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1595 U$$3946/B1 VGND VGND VPWR VPWR U$$384/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_66_1 dadda_fa_5_66_1/A dadda_fa_5_66_1/B dadda_fa_5_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_67_0/B dadda_fa_7_66_0/A sky130_fd_sc_hd__fa_2
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_59_0 dadda_fa_5_59_0/A dadda_fa_5_59_0/B dadda_fa_5_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_60_0/A dadda_fa_6_59_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_141_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_58_8 dadda_fa_1_58_8/A dadda_fa_1_58_8/B dadda_fa_1_58_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_59_3/A dadda_fa_3_58_0/A sky130_fd_sc_hd__fa_2
XFILLER_82_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_105_0 U$$2876/Y U$$3010/X U$$3143/X VGND VGND VPWR VPWR dadda_fa_3_106_3/A
+ dadda_fa_3_105_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_165_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2080 U$$2080/A U$$2094/B VGND VGND VPWR VPWR U$$2080/X sky130_fd_sc_hd__xor2_1
XFILLER_210_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2091 U$$4009/A1 U$$2091/A2 U$$860/A1 U$$2091/B2 VGND VGND VPWR VPWR U$$2092/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1390 U$$1799/B1 U$$1422/A2 U$$1666/A1 U$$1422/B2 VGND VGND VPWR VPWR U$$1391/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_496 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_91_2 U$$2716/X U$$2849/X U$$2982/X VGND VGND VPWR VPWR dadda_fa_2_92_5/A
+ dadda_fa_3_91_0/A sky130_fd_sc_hd__fa_2
XFILLER_191_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_84_1 U$$1771/X U$$1904/X U$$2037/X VGND VGND VPWR VPWR dadda_fa_2_85_2/B
+ dadda_fa_2_84_4/B sky130_fd_sc_hd__fa_1
XFILLER_104_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_61_0 dadda_fa_4_61_0/A dadda_fa_4_61_0/B dadda_fa_4_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/A dadda_fa_5_61_1/A sky130_fd_sc_hd__fa_1
XFILLER_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_77_0 U$$1358/X U$$1491/X U$$1624/X VGND VGND VPWR VPWR dadda_fa_2_78_0/B
+ dadda_fa_2_77_3/B sky130_fd_sc_hd__fa_1
XTAP_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_2_104_2 U$$3540/X U$$3673/X VGND VGND VPWR VPWR dadda_fa_3_105_3/B dadda_fa_4_104_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3709 U$$832/A1 U$$3793/A2 U$$3846/B1 U$$3793/B2 VGND VGND VPWR VPWR U$$3710/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1006 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_328 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_373_ _373_/CLK _373_/D VGND VGND VPWR VPWR _373_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_207_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4399_1776 VGND VGND VPWR VPWR U$$4399_1776/HI U$$4399/B sky130_fd_sc_hd__conb_1
XFILLER_182_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_99_1 dadda_fa_3_99_1/A dadda_fa_3_99_1/B dadda_fa_3_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_0/CIN dadda_fa_4_99_2/A sky130_fd_sc_hd__fa_1
XFILLER_127_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_76_0 dadda_fa_6_76_0/A dadda_fa_6_76_0/B dadda_fa_6_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_77_0/B dadda_fa_7_76_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_859 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$470 U$$470/A U$$474/B VGND VGND VPWR VPWR U$$470/X sky130_fd_sc_hd__xor2_1
XU$$481 U$$616/B1 U$$483/A2 U$$757/A1 U$$483/B2 VGND VGND VPWR VPWR U$$482/A sky130_fd_sc_hd__a22o_1
XFILLER_205_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$492 U$$492/A U$$492/B VGND VGND VPWR VPWR U$$492/X sky130_fd_sc_hd__xor2_1
XFILLER_149_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_94_0 U$$2722/X U$$2855/X U$$2988/X VGND VGND VPWR VPWR dadda_fa_3_95_0/B
+ dadda_fa_3_94_2/B sky130_fd_sc_hd__fa_1
XFILLER_133_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1370 U$$2543/B VGND VGND VPWR VPWR U$$2525/B sky130_fd_sc_hd__buf_6
XFILLER_132_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1381 U$$796/B VGND VGND VPWR VPWR U$$750/B sky130_fd_sc_hd__buf_6
XFILLER_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1392 input29/X VGND VGND VPWR VPWR U$$2466/A sky130_fd_sc_hd__buf_6
XFILLER_114_886 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_70_7 dadda_fa_1_70_7/A dadda_fa_1_70_7/B dadda_fa_1_70_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_2/CIN dadda_fa_2_70_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_6 dadda_fa_1_63_6/A dadda_fa_1_63_6/B dadda_fa_1_63_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_2/B dadda_fa_2_63_5/B sky130_fd_sc_hd__fa_1
XFILLER_80_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_56_5 U$$3178/X U$$3311/X U$$3444/X VGND VGND VPWR VPWR dadda_fa_2_57_2/A
+ dadda_fa_2_56_5/A sky130_fd_sc_hd__fa_1
XFILLER_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_49_4 U$$1701/X U$$1834/X U$$1967/X VGND VGND VPWR VPWR dadda_fa_2_50_2/A
+ dadda_fa_2_49_5/A sky130_fd_sc_hd__fa_1
XFILLER_55_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_19_2 dadda_fa_4_19_2/A dadda_fa_4_19_2/B dadda_ha_3_19_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_20_0/CIN dadda_fa_5_19_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_202_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_93_0 dadda_fa_7_93_0/A dadda_fa_7_93_0/B dadda_fa_7_93_0/CIN VGND VGND
+ VPWR VPWR _390_/D _261_/D sky130_fd_sc_hd__fa_2
XFILLER_13_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4207 U$$4207/A U$$4211/B VGND VGND VPWR VPWR U$$4207/X sky130_fd_sc_hd__xor2_1
XFILLER_133_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4218 input110/X U$$4240/A2 input111/X U$$4240/B2 VGND VGND VPWR VPWR U$$4219/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4229 U$$4229/A U$$4239/B VGND VGND VPWR VPWR U$$4229/X sky130_fd_sc_hd__xor2_1
XFILLER_93_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3506 U$$3506/A U$$3510/B VGND VGND VPWR VPWR U$$3506/X sky130_fd_sc_hd__xor2_1
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3517 U$$3517/A1 U$$3517/A2 U$$4478/A1 U$$3517/B2 VGND VGND VPWR VPWR U$$3518/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3528 U$$3528/A U$$3528/B VGND VGND VPWR VPWR U$$3528/X sky130_fd_sc_hd__xor2_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3539 U$$3813/A1 U$$3549/A2 U$$116/A1 U$$3549/B2 VGND VGND VPWR VPWR U$$3540/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2805 U$$2805/A U$$2825/B VGND VGND VPWR VPWR U$$2805/X sky130_fd_sc_hd__xor2_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2816 U$$2951/B1 U$$2828/A2 U$$4323/B1 U$$2828/B2 VGND VGND VPWR VPWR U$$2817/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2827 U$$2827/A U$$2845/B VGND VGND VPWR VPWR U$$2827/X sky130_fd_sc_hd__xor2_1
XU$$2838 U$$2975/A1 U$$2744/X U$$2975/B1 U$$2745/X VGND VGND VPWR VPWR U$$2839/A sky130_fd_sc_hd__a22o_1
XANTENNA_121 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 _237_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2849 U$$2849/A U$$2876/A VGND VGND VPWR VPWR U$$2849/X sky130_fd_sc_hd__xor2_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_21_2 U$$847/X U$$980/X U$$1113/X VGND VGND VPWR VPWR dadda_fa_4_22_1/A
+ dadda_fa_4_21_2/B sky130_fd_sc_hd__fa_1
XANTENNA_143 U$$1877/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 U$$2828/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_165 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_176 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_187 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_198 _199_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_356_ _359_/CLK _356_/D VGND VGND VPWR VPWR _356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_287_ _417_/CLK _287_/D VGND VGND VPWR VPWR _287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_73_5 dadda_fa_2_73_5/A dadda_fa_2_73_5/B dadda_fa_2_73_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_74_2/A dadda_fa_4_73_0/A sky130_fd_sc_hd__fa_1
XFILLER_25_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_66_4 dadda_fa_2_66_4/A dadda_fa_2_66_4/B dadda_fa_2_66_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_1/CIN dadda_fa_3_66_3/CIN sky130_fd_sc_hd__fa_2
XFILLER_96_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_59_3 dadda_fa_2_59_3/A dadda_fa_2_59_3/B dadda_fa_2_59_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/B dadda_fa_3_59_3/B sky130_fd_sc_hd__fa_1
XFILLER_110_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 a[13] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__buf_4
XFILLER_65_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1095 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_29_1 dadda_fa_5_29_1/A dadda_fa_5_29_1/B dadda_fa_5_29_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_30_0/B dadda_fa_7_29_0/A sky130_fd_sc_hd__fa_1
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_934 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$3 _299_/Q _171_/Q VGND VGND VPWR VPWR final_adder.U$$3/COUT final_adder.U$$3/SUM
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_5_103_1 dadda_fa_5_103_1/A dadda_fa_5_103_1/B dadda_fa_5_103_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_104_0/B dadda_fa_7_103_0/A sky130_fd_sc_hd__fa_2
XFILLER_173_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput320 output320/A VGND VGND VPWR VPWR o[41] sky130_fd_sc_hd__buf_2
XFILLER_161_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput331 output331/A VGND VGND VPWR VPWR o[51] sky130_fd_sc_hd__buf_2
XFILLER_126_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput342 output342/A VGND VGND VPWR VPWR o[61] sky130_fd_sc_hd__buf_2
Xoutput353 output353/A VGND VGND VPWR VPWR o[71] sky130_fd_sc_hd__buf_2
Xoutput364 output364/A VGND VGND VPWR VPWR o[81] sky130_fd_sc_hd__buf_2
Xoutput375 output375/A VGND VGND VPWR VPWR o[91] sky130_fd_sc_hd__buf_2
XFILLER_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_61_3 U$$3188/X U$$3321/X U$$3454/X VGND VGND VPWR VPWR dadda_fa_2_62_1/B
+ dadda_fa_2_61_4/B sky130_fd_sc_hd__fa_1
XFILLER_101_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_2 U$$1578/X U$$1711/X U$$1844/X VGND VGND VPWR VPWR dadda_fa_2_55_1/A
+ dadda_fa_2_54_4/A sky130_fd_sc_hd__fa_1
XFILLER_56_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_31_1 dadda_fa_4_31_1/A dadda_fa_4_31_1/B dadda_fa_4_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/B dadda_fa_5_31_1/B sky130_fd_sc_hd__fa_1
XFILLER_132_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_47_1 U$$500/X U$$633/X U$$766/X VGND VGND VPWR VPWR dadda_fa_2_48_1/CIN
+ dadda_fa_2_47_4/B sky130_fd_sc_hd__fa_1
XFILLER_71_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_24_0 dadda_fa_4_24_0/A dadda_fa_4_24_0/B dadda_fa_4_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/A dadda_fa_5_24_1/A sky130_fd_sc_hd__fa_1
XFILLER_167_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_210_ _211_/CLK _210_/D VGND VGND VPWR VPWR _210_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_196_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_274 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_76_3 dadda_fa_3_76_3/A dadda_fa_3_76_3/B dadda_fa_3_76_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_77_1/B dadda_fa_4_76_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_111_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_69_2 dadda_fa_3_69_2/A dadda_fa_3_69_2/B dadda_fa_3_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_1/A dadda_fa_4_69_2/B sky130_fd_sc_hd__fa_1
XFILLER_78_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4004 U$$4004/A U$$4036/B VGND VGND VPWR VPWR U$$4004/X sky130_fd_sc_hd__xor2_1
XFILLER_76_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4015 input73/X U$$4079/A2 U$$4015/B1 U$$4079/B2 VGND VGND VPWR VPWR U$$4016/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4026 U$$4026/A U$$4044/B VGND VGND VPWR VPWR U$$4026/X sky130_fd_sc_hd__xor2_1
XU$$4037 U$$4309/B1 U$$3977/X U$$4176/A1 U$$3978/X VGND VGND VPWR VPWR U$$4038/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_39_0 dadda_fa_6_39_0/A dadda_fa_6_39_0/B dadda_fa_6_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_40_0/B dadda_fa_7_39_0/CIN sky130_fd_sc_hd__fa_1
XU$$3303 U$$3303/A U$$3395/B VGND VGND VPWR VPWR U$$3303/X sky130_fd_sc_hd__xor2_1
XU$$4048 U$$4048/A U$$4100/B VGND VGND VPWR VPWR U$$4048/X sky130_fd_sc_hd__xor2_1
XFILLER_76_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4059 U$$4333/A1 U$$4077/A2 U$$4333/B1 U$$4077/B2 VGND VGND VPWR VPWR U$$4060/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3314 U$$3451/A1 U$$3320/A2 U$$711/B1 U$$3320/B2 VGND VGND VPWR VPWR U$$3315/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3325 U$$3325/A U$$3349/B VGND VGND VPWR VPWR U$$3325/X sky130_fd_sc_hd__xor2_1
XFILLER_47_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3336 U$$4432/A1 U$$3292/X U$$4434/A1 U$$3293/X VGND VGND VPWR VPWR U$$3337/A sky130_fd_sc_hd__a22o_1
XFILLER_207_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2602 U$$2602/A VGND VGND VPWR VPWR U$$2602/Y sky130_fd_sc_hd__inv_1
XU$$3347 U$$3347/A U$$3349/B VGND VGND VPWR VPWR U$$3347/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2613 U$$3296/B1 U$$2625/A2 U$$3026/A1 U$$2625/B2 VGND VGND VPWR VPWR U$$2614/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3358 U$$4178/B1 U$$3378/A2 U$$4045/A1 U$$3378/B2 VGND VGND VPWR VPWR U$$3359/A
+ sky130_fd_sc_hd__a22o_1
XU$$3369 U$$3369/A U$$3375/B VGND VGND VPWR VPWR U$$3369/X sky130_fd_sc_hd__xor2_1
XU$$2624 U$$2624/A U$$2624/B VGND VGND VPWR VPWR U$$2624/X sky130_fd_sc_hd__xor2_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2635 U$$3183/A1 U$$2653/A2 U$$3183/B1 U$$2653/B2 VGND VGND VPWR VPWR U$$2636/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1901 U$$2312/A1 U$$1913/A2 U$$2312/B1 U$$1903/B2 VGND VGND VPWR VPWR U$$1902/A
+ sky130_fd_sc_hd__a22o_1
XU$$2646 U$$2646/A U$$2650/B VGND VGND VPWR VPWR U$$2646/X sky130_fd_sc_hd__xor2_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1912 U$$1912/A U$$1912/B VGND VGND VPWR VPWR U$$1912/X sky130_fd_sc_hd__xor2_1
XU$$2657 U$$874/B1 U$$2683/A2 U$$330/A1 U$$2683/B2 VGND VGND VPWR VPWR U$$2658/A sky130_fd_sc_hd__a22o_1
XFILLER_62_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2668 U$$2668/A U$$2710/B VGND VGND VPWR VPWR U$$2668/X sky130_fd_sc_hd__xor2_1
XU$$1923 U$$1921/B input20/X input21/X U$$1918/Y VGND VGND VPWR VPWR U$$1923/X sky130_fd_sc_hd__a22o_2
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2679 U$$3499/B1 U$$2691/A2 U$$2955/A1 U$$2691/B2 VGND VGND VPWR VPWR U$$2680/A
+ sky130_fd_sc_hd__a22o_1
XU$$1934 U$$2206/B1 U$$1970/A2 U$$3032/A1 U$$1970/B2 VGND VGND VPWR VPWR U$$1935/A
+ sky130_fd_sc_hd__a22o_1
XU$$1945 U$$1945/A U$$2009/B VGND VGND VPWR VPWR U$$1945/X sky130_fd_sc_hd__xor2_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1956 U$$860/A1 U$$2040/A2 U$$860/B1 U$$2040/B2 VGND VGND VPWR VPWR U$$1957/A sky130_fd_sc_hd__a22o_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1967 U$$1967/A U$$1971/B VGND VGND VPWR VPWR U$$1967/X sky130_fd_sc_hd__xor2_1
XU$$1978 U$$2113/B1 U$$2016/A2 U$$3348/B1 U$$2016/B2 VGND VGND VPWR VPWR U$$1979/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_408_ _408_/CLK _408_/D VGND VGND VPWR VPWR _408_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1989 U$$1989/A U$$1991/B VGND VGND VPWR VPWR U$$1989/X sky130_fd_sc_hd__xor2_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_339_ _342_/CLK _339_/D VGND VGND VPWR VPWR _339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_414 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_71_2 dadda_fa_2_71_2/A dadda_fa_2_71_2/B dadda_fa_2_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/A dadda_fa_3_71_3/A sky130_fd_sc_hd__fa_1
XFILLER_29_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_64_1 dadda_fa_2_64_1/A dadda_fa_2_64_1/B dadda_fa_2_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_0/CIN dadda_fa_3_64_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater801 U$$2435/B2 VGND VGND VPWR VPWR U$$2417/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$608 final_adder.U$$616/B final_adder.U$$608/B VGND VGND VPWR VPWR
+ final_adder.U$$712/A sky130_fd_sc_hd__and2_1
Xrepeater812 U$$2197/X VGND VGND VPWR VPWR U$$2316/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_110_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$619 final_adder.U$$610/A final_adder.U$$503/X final_adder.U$$495/X
+ VGND VGND VPWR VPWR final_adder.U$$619/X sky130_fd_sc_hd__a21o_2
Xdadda_fa_5_41_0 dadda_fa_5_41_0/A dadda_fa_5_41_0/B dadda_fa_5_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_42_0/A dadda_fa_6_41_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater823 U$$1990/B2 VGND VGND VPWR VPWR U$$1970/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_57_0 dadda_fa_2_57_0/A dadda_fa_2_57_0/B dadda_fa_2_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_0/B dadda_fa_3_57_2/B sky130_fd_sc_hd__fa_1
Xrepeater834 U$$1903/B2 VGND VGND VPWR VPWR U$$1877/B2 sky130_fd_sc_hd__buf_8
XFILLER_38_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater845 U$$1770/B2 VGND VGND VPWR VPWR U$$1746/B2 sky130_fd_sc_hd__buf_8
XFILLER_84_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater856 U$$175/B2 VGND VGND VPWR VPWR U$$165/B2 sky130_fd_sc_hd__buf_2
Xrepeater867 U$$1462/B2 VGND VGND VPWR VPWR U$$1434/B2 sky130_fd_sc_hd__buf_6
Xrepeater878 U$$1238/X VGND VGND VPWR VPWR U$$1337/B2 sky130_fd_sc_hd__buf_6
XFILLER_37_431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$30 U$$30/A1 U$$50/A2 U$$32/A1 U$$50/B2 VGND VGND VPWR VPWR U$$31/A sky130_fd_sc_hd__a22o_1
Xrepeater889 U$$50/B2 VGND VGND VPWR VPWR U$$42/B2 sky130_fd_sc_hd__buf_2
XU$$41 U$$41/A U$$43/B VGND VGND VPWR VPWR U$$41/X sky130_fd_sc_hd__xor2_1
XFILLER_37_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$52 U$$52/A1 U$$80/A2 U$$52/B1 U$$80/B2 VGND VGND VPWR VPWR U$$53/A sky130_fd_sc_hd__a22o_1
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$63 U$$63/A U$$85/B VGND VGND VPWR VPWR U$$63/X sky130_fd_sc_hd__xor2_1
XFILLER_37_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_935 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$74 U$$74/A1 U$$80/A2 U$$76/A1 U$$80/B2 VGND VGND VPWR VPWR U$$75/A sky130_fd_sc_hd__a22o_1
XU$$85 U$$85/A U$$85/B VGND VGND VPWR VPWR U$$85/X sky130_fd_sc_hd__xor2_1
XU$$3870 U$$4418/A1 U$$3902/A2 U$$4420/A1 U$$3902/B2 VGND VGND VPWR VPWR U$$3871/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_198_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$96 U$$96/A1 U$$98/A2 U$$98/A1 U$$98/B2 VGND VGND VPWR VPWR U$$97/A sky130_fd_sc_hd__a22o_1
XU$$3881 U$$3881/A U$$3971/B VGND VGND VPWR VPWR U$$3881/X sky130_fd_sc_hd__xor2_1
XFILLER_198_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3892 U$$4029/A1 U$$3970/A2 input82/X U$$3970/B2 VGND VGND VPWR VPWR U$$3893/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_607 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_10 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_21 _336_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_32 _339_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_43 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_634 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_54 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_65 _342_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_76 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_807 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_87 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_197_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_98 _346_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_86_2 dadda_fa_4_86_2/A dadda_fa_4_86_2/B dadda_fa_4_86_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_87_0/CIN dadda_fa_5_86_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_79_1 dadda_fa_4_79_1/A dadda_fa_4_79_1/B dadda_fa_4_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/B dadda_fa_5_79_1/B sky130_fd_sc_hd__fa_1
XFILLER_47_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_56_0 dadda_fa_7_56_0/A dadda_fa_7_56_0/B dadda_fa_7_56_0/CIN VGND VGND
+ VPWR VPWR _353_/D _224_/D sky130_fd_sc_hd__fa_1
XFILLER_134_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_718 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1208 U$$932/B1 U$$1100/X U$$799/A1 U$$1101/X VGND VGND VPWR VPWR U$$1209/A sky130_fd_sc_hd__a22o_1
XU$$1219 U$$1219/A U$$1232/A VGND VGND VPWR VPWR U$$1219/X sky130_fd_sc_hd__xor2_1
XFILLER_204_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1013 final_adder.U$$242/A final_adder.U$$623/X final_adder.U$$243/A2
+ VGND VGND VPWR VPWR final_adder.U$$1037/B sky130_fd_sc_hd__a21o_1
XFILLER_89_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1024 final_adder.U$$0/SUM final_adder.U$$1024/B VGND VGND VPWR VPWR
+ output257/A sky130_fd_sc_hd__xor2_1
XFILLER_8_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$1035 final_adder.U$$244/B final_adder.U$$1035/B VGND VGND VPWR VPWR
+ output279/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1046 final_adder.U$$232/A final_adder.U$$733/X VGND VGND VPWR VPWR
+ output299/A sky130_fd_sc_hd__xor2_1
XFILLER_137_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1057 final_adder.U$$222/B final_adder.U$$993/X VGND VGND VPWR VPWR
+ output311/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1068 final_adder.U$$210/A final_adder.U$$823/X VGND VGND VPWR VPWR
+ output323/A sky130_fd_sc_hd__xor2_1
XFILLER_165_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$1079 final_adder.U$$200/B final_adder.U$$971/X VGND VGND VPWR VPWR
+ output335/A sky130_fd_sc_hd__xor2_1
XFILLER_109_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_81_1 dadda_fa_3_81_1/A dadda_fa_3_81_1/B dadda_fa_3_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_0/CIN dadda_fa_4_81_2/A sky130_fd_sc_hd__fa_1
XFILLER_178_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_74_0 dadda_fa_3_74_0/A dadda_fa_3_74_0/B dadda_fa_3_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_0/B dadda_fa_4_74_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_106_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3100 U$$3235/B1 U$$3108/A2 U$$3376/A1 U$$3108/B2 VGND VGND VPWR VPWR U$$3101/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3111 U$$3111/A U$$3151/A VGND VGND VPWR VPWR U$$3111/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_110_1 dadda_fa_4_110_1/A dadda_fa_4_110_1/B dadda_fa_4_110_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_111_0/B dadda_fa_5_110_1/B sky130_fd_sc_hd__fa_1
XU$$3122 U$$517/B1 U$$3132/A2 U$$384/A1 U$$3132/B2 VGND VGND VPWR VPWR U$$3123/A sky130_fd_sc_hd__a22o_1
XU$$3133 U$$3133/A U$$3133/B VGND VGND VPWR VPWR U$$3133/X sky130_fd_sc_hd__xor2_1
XU$$3144 input122/X U$$3148/A2 U$$3281/B1 U$$3148/B2 VGND VGND VPWR VPWR U$$3145/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2410 U$$2410/A U$$2426/B VGND VGND VPWR VPWR U$$2410/X sky130_fd_sc_hd__xor2_1
XU$$3155 U$$3153/Y input41/X U$$3151/A U$$3154/X U$$3151/Y VGND VGND VPWR VPWR U$$3155/X
+ sky130_fd_sc_hd__a32o_4
Xdadda_fa_2_36_5 input186/X dadda_fa_2_36_5/B dadda_fa_2_36_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_37_2/A dadda_fa_4_36_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_103_0 dadda_fa_4_103_0/A dadda_fa_4_103_0/B dadda_fa_4_103_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/A dadda_fa_5_103_1/A sky130_fd_sc_hd__fa_1
XU$$3166 U$$3166/A U$$3188/B VGND VGND VPWR VPWR U$$3166/X sky130_fd_sc_hd__xor2_1
XU$$2421 U$$366/A1 U$$2459/A2 U$$3245/A1 U$$2459/B2 VGND VGND VPWR VPWR U$$2422/A
+ sky130_fd_sc_hd__a22o_1
XU$$3177 U$$3451/A1 U$$3263/A2 input66/X U$$3263/B2 VGND VGND VPWR VPWR U$$3178/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2432 U$$2432/A U$$2466/A VGND VGND VPWR VPWR U$$2432/X sky130_fd_sc_hd__xor2_1
XU$$2443 U$$936/A1 U$$2333/X U$$936/B1 U$$2334/X VGND VGND VPWR VPWR U$$2444/A sky130_fd_sc_hd__a22o_1
XFILLER_46_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3188 U$$3188/A U$$3188/B VGND VGND VPWR VPWR U$$3188/X sky130_fd_sc_hd__xor2_1
XU$$2454 U$$2454/A U$$2454/B VGND VGND VPWR VPWR U$$2454/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3199 U$$4432/A1 U$$3241/A2 U$$4434/A1 U$$3241/B2 VGND VGND VPWR VPWR U$$3200/A
+ sky130_fd_sc_hd__a22o_1
XU$$1720 U$$2951/B1 U$$1750/A2 U$$78/A1 U$$1750/B2 VGND VGND VPWR VPWR U$$1721/A sky130_fd_sc_hd__a22o_1
XU$$2465 U$$2465/A VGND VGND VPWR VPWR U$$2465/Y sky130_fd_sc_hd__inv_1
XFILLER_146_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1731 U$$1731/A U$$1739/B VGND VGND VPWR VPWR U$$1731/X sky130_fd_sc_hd__xor2_1
XU$$2476 U$$3296/B1 U$$2524/A2 U$$3026/A1 U$$2524/B2 VGND VGND VPWR VPWR U$$2477/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2487 U$$2487/A U$$2491/B VGND VGND VPWR VPWR U$$2487/X sky130_fd_sc_hd__xor2_1
XU$$1742 U$$2016/A1 U$$1770/A2 U$$2701/B1 U$$1770/B2 VGND VGND VPWR VPWR U$$1743/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1753 U$$1753/A U$$1765/B VGND VGND VPWR VPWR U$$1753/X sky130_fd_sc_hd__xor2_1
XFILLER_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2498 U$$3183/A1 U$$2542/A2 U$$3183/B1 U$$2542/B2 VGND VGND VPWR VPWR U$$2499/A
+ sky130_fd_sc_hd__a22o_1
XU$$1764 U$$2449/A1 U$$1764/A2 U$$1764/B1 U$$1764/B2 VGND VGND VPWR VPWR U$$1765/A
+ sky130_fd_sc_hd__a22o_1
XU$$1775 U$$1775/A U$$1779/B VGND VGND VPWR VPWR U$$1775/X sky130_fd_sc_hd__xor2_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1786 U$$1784/B input18/X input19/X U$$1781/Y VGND VGND VPWR VPWR U$$1786/X sky130_fd_sc_hd__a22o_4
XFILLER_175_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1797 U$$1932/B1 U$$1831/A2 U$$1799/A1 U$$1831/B2 VGND VGND VPWR VPWR U$$1798/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_96_1 dadda_fa_5_96_1/A dadda_fa_5_96_1/B dadda_fa_5_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_97_0/B dadda_fa_7_96_0/A sky130_fd_sc_hd__fa_1
XFILLER_135_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 a[36] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 a[46] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 a[56] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput63 a[8] VGND VGND VPWR VPWR U$$549/A sky130_fd_sc_hd__buf_2
XFILLER_200_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_892 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_89_0 dadda_fa_5_89_0/A dadda_fa_5_89_0/B dadda_fa_5_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_90_0/A dadda_fa_6_89_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_115_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput74 b[18] VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__buf_8
XFILLER_7_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput85 b[28] VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__buf_8
XFILLER_155_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput96 b[38] VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__buf_6
XFILLER_192_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$405 final_adder.U$$404/B final_adder.U$$283/X final_adder.U$$279/X
+ VGND VGND VPWR VPWR final_adder.U$$405/X sky130_fd_sc_hd__a21o_1
XFILLER_85_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$416 final_adder.U$$420/B final_adder.U$$416/B VGND VGND VPWR VPWR
+ final_adder.U$$540/B sky130_fd_sc_hd__and2_1
Xrepeater620 U$$1462/A2 VGND VGND VPWR VPWR U$$1434/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$427 final_adder.U$$426/B final_adder.U$$305/X final_adder.U$$301/X
+ VGND VGND VPWR VPWR final_adder.U$$427/X sky130_fd_sc_hd__a21o_1
Xrepeater631 U$$1237/X VGND VGND VPWR VPWR U$$1367/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$438 final_adder.U$$442/B final_adder.U$$438/B VGND VGND VPWR VPWR
+ final_adder.U$$562/B sky130_fd_sc_hd__and2_1
XTAP_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater642 U$$1057/B2 VGND VGND VPWR VPWR U$$979/B2 sky130_fd_sc_hd__buf_4
XFILLER_123_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$449 final_adder.U$$448/B final_adder.U$$327/X final_adder.U$$323/X
+ VGND VGND VPWR VPWR final_adder.U$$449/X sky130_fd_sc_hd__a21o_1
Xrepeater653 U$$938/B2 VGND VGND VPWR VPWR U$$950/B2 sky130_fd_sc_hd__buf_8
XFILLER_84_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater664 U$$636/B2 VGND VGND VPWR VPWR U$$606/B2 sky130_fd_sc_hd__buf_4
Xrepeater675 U$$4369/B2 VGND VGND VPWR VPWR U$$4361/B2 sky130_fd_sc_hd__buf_4
XFILLER_44_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater686 U$$4164/B2 VGND VGND VPWR VPWR U$$4144/B2 sky130_fd_sc_hd__buf_4
Xrepeater697 U$$4103/B2 VGND VGND VPWR VPWR U$$4079/B2 sky130_fd_sc_hd__buf_4
XU$$4386_1767 VGND VGND VPWR VPWR U$$4386_1767/HI U$$4386/A sky130_fd_sc_hd__conb_1
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4390 U$$4390/A1 U$$4388/X U$$4392/A1 U$$4432/B2 VGND VGND VPWR VPWR U$$4391/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_91_0 dadda_fa_4_91_0/A dadda_fa_4_91_0/B ANTENNA_0/DIODE VGND VGND VPWR
+ VPWR dadda_fa_5_92_0/A dadda_fa_5_91_1/A sky130_fd_sc_hd__fa_1
XFILLER_140_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_583 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_105_2 U$$4473/X input135/X dadda_fa_3_105_2/CIN VGND VGND VPWR VPWR dadda_fa_4_106_1/A
+ dadda_fa_4_105_2/B sky130_fd_sc_hd__fa_1
XFILLER_107_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_119_0 dadda_fa_6_119_0/A dadda_fa_6_119_0/B dadda_fa_6_119_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_120_0/B dadda_fa_7_119_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$961 final_adder.U$$190/A final_adder.U$$803/X final_adder.U$$961/B1
+ VGND VGND VPWR VPWR final_adder.U$$961/X sky130_fd_sc_hd__a21o_1
XU$$800 U$$800/A U$$808/B VGND VGND VPWR VPWR U$$800/X sky130_fd_sc_hd__xor2_1
XTAP_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$811 U$$811/A1 U$$689/X U$$950/A1 U$$690/X VGND VGND VPWR VPWR U$$812/A sky130_fd_sc_hd__a22o_1
XFILLER_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$983 final_adder.U$$212/A final_adder.U$$825/X final_adder.U$$983/B1
+ VGND VGND VPWR VPWR final_adder.U$$983/X sky130_fd_sc_hd__a21o_1
XU$$822 input3/X VGND VGND VPWR VPWR U$$822/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_3_39_3 dadda_fa_3_39_3/A dadda_fa_3_39_3/B dadda_fa_3_39_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_40_1/B dadda_fa_4_39_2/CIN sky130_fd_sc_hd__fa_1
XU$$833 U$$833/A U$$847/B VGND VGND VPWR VPWR U$$833/X sky130_fd_sc_hd__xor2_1
XFILLER_17_935 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$844 U$$981/A1 U$$906/A2 U$$983/A1 U$$906/B2 VGND VGND VPWR VPWR U$$845/A sky130_fd_sc_hd__a22o_1
XFILLER_189_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$855 U$$855/A U$$877/B VGND VGND VPWR VPWR U$$855/X sky130_fd_sc_hd__xor2_1
XU$$866 U$$866/A1 U$$882/A2 U$$46/A1 U$$882/B2 VGND VGND VPWR VPWR U$$867/A sky130_fd_sc_hd__a22o_1
XU$$1005 U$$46/A1 U$$999/A2 U$$48/A1 U$$999/B2 VGND VGND VPWR VPWR U$$1006/A sky130_fd_sc_hd__a22o_1
XU$$1016 U$$1016/A U$$998/B VGND VGND VPWR VPWR U$$1016/X sky130_fd_sc_hd__xor2_1
XU$$877 U$$877/A U$$877/B VGND VGND VPWR VPWR U$$877/X sky130_fd_sc_hd__xor2_1
XU$$1027 U$$890/A1 U$$1083/A2 U$$892/A1 U$$1083/B2 VGND VGND VPWR VPWR U$$1028/A sky130_fd_sc_hd__a22o_1
XU$$888 U$$888/A1 U$$892/A2 U$$890/A1 U$$892/B2 VGND VGND VPWR VPWR U$$889/A sky130_fd_sc_hd__a22o_1
XU$$899 U$$899/A U$$951/B VGND VGND VPWR VPWR U$$899/X sky130_fd_sc_hd__xor2_1
XU$$1038 U$$1038/A U$$980/B VGND VGND VPWR VPWR U$$1038/X sky130_fd_sc_hd__xor2_1
XFILLER_189_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1049 U$$773/B1 U$$965/A2 U$$640/A1 U$$965/B2 VGND VGND VPWR VPWR U$$1050/A sky130_fd_sc_hd__a22o_1
XFILLER_204_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1700 input101/X VGND VGND VPWR VPWR U$$3517/A1 sky130_fd_sc_hd__buf_4
XFILLER_32_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_927 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_ha_2_28_3 U$$1260/X U$$1393/X VGND VGND VPWR VPWR dadda_fa_3_29_2/CIN dadda_fa_4_28_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_6_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1036 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_41_3 U$$2749/X input192/X dadda_fa_2_41_3/CIN VGND VGND VPWR VPWR dadda_fa_3_42_1/B
+ dadda_fa_3_41_3/B sky130_fd_sc_hd__fa_1
XFILLER_81_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_34_2 U$$1139/X U$$1272/X U$$1405/X VGND VGND VPWR VPWR dadda_fa_3_35_1/A
+ dadda_fa_3_34_3/A sky130_fd_sc_hd__fa_1
XFILLER_207_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_11_1 dadda_fa_5_11_1/A dadda_fa_5_11_1/B dadda_ha_4_11_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_12_0/B dadda_fa_7_11_0/A sky130_fd_sc_hd__fa_1
XU$$2240 U$$3882/B1 U$$2284/A2 U$$3749/A1 U$$2284/B2 VGND VGND VPWR VPWR U$$2241/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2251 U$$2251/A U$$2253/B VGND VGND VPWR VPWR U$$2251/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_27_1 U$$460/X U$$593/X U$$726/X VGND VGND VPWR VPWR dadda_fa_3_28_2/B
+ dadda_fa_3_27_3/CIN sky130_fd_sc_hd__fa_1
XU$$2262 U$$892/A1 U$$2308/A2 U$$894/A1 U$$2308/B2 VGND VGND VPWR VPWR U$$2263/A sky130_fd_sc_hd__a22o_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2273 U$$2273/A U$$2273/B VGND VGND VPWR VPWR U$$2273/X sky130_fd_sc_hd__xor2_1
XU$$2284 U$$914/A1 U$$2284/A2 U$$914/B1 U$$2284/B2 VGND VGND VPWR VPWR U$$2285/A sky130_fd_sc_hd__a22o_1
XFILLER_195_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1550 U$$1550/A U$$1558/B VGND VGND VPWR VPWR U$$1550/X sky130_fd_sc_hd__xor2_1
XU$$2295 U$$2295/A U$$2317/B VGND VGND VPWR VPWR U$$2295/X sky130_fd_sc_hd__xor2_1
XFILLER_167_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1561 U$$874/B1 U$$1591/A2 U$$330/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1562/A sky130_fd_sc_hd__a22o_1
XU$$1572 U$$1572/A U$$1574/B VGND VGND VPWR VPWR U$$1572/X sky130_fd_sc_hd__xor2_1
XFILLER_195_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1583 U$$2951/B1 U$$1621/A2 U$$4323/B1 U$$1621/B2 VGND VGND VPWR VPWR U$$1584/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1594 U$$1594/A U$$1608/B VGND VGND VPWR VPWR U$$1594/X sky130_fd_sc_hd__xor2_1
XFILLER_163_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_79_4 U$$2692/X U$$2825/X U$$2958/X VGND VGND VPWR VPWR dadda_fa_2_80_1/CIN
+ dadda_fa_2_79_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$202 final_adder.U$$202/A final_adder.U$$202/B VGND VGND VPWR VPWR
+ final_adder.U$$330/B sky130_fd_sc_hd__and2_1
XTAP_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$213 final_adder.U$$212/B final_adder.U$$983/B1 final_adder.U$$213/B1
+ VGND VGND VPWR VPWR final_adder.U$$213/X sky130_fd_sc_hd__a21o_1
XTAP_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$224 final_adder.U$$224/A final_adder.U$$224/B VGND VGND VPWR VPWR
+ final_adder.U$$352/B sky130_fd_sc_hd__and2_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_49_2 dadda_fa_4_49_2/A dadda_fa_4_49_2/B dadda_fa_4_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_50_0/CIN dadda_fa_5_49_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_111_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$235 final_adder.U$$234/B final_adder.U$$235/A2 final_adder.U$$235/B1
+ VGND VGND VPWR VPWR final_adder.U$$235/X sky130_fd_sc_hd__a21o_1
XTAP_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$246 final_adder.U$$8/SUM final_adder.U$$9/SUM VGND VGND VPWR VPWR
+ final_adder.U$$374/B sky130_fd_sc_hd__and2_1
Xrepeater450 U$$4103/A2 VGND VGND VPWR VPWR U$$4079/A2 sky130_fd_sc_hd__buf_4
XTAP_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater461 U$$3968/A2 VGND VGND VPWR VPWR U$$3966/A2 sky130_fd_sc_hd__buf_8
Xfinal_adder.U$$268 final_adder.U$$270/B final_adder.U$$268/B VGND VGND VPWR VPWR
+ final_adder.U$$394/B sky130_fd_sc_hd__and2_1
XTAP_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater472 U$$3644/A2 VGND VGND VPWR VPWR U$$3612/A2 sky130_fd_sc_hd__clkbuf_8
XU$$107 U$$107/A U$$111/B VGND VGND VPWR VPWR U$$107/X sky130_fd_sc_hd__xor2_1
XFILLER_211_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$279 final_adder.U$$278/B final_adder.U$$153/X final_adder.U$$151/X
+ VGND VGND VPWR VPWR final_adder.U$$279/X sky130_fd_sc_hd__a21o_1
XU$$118 U$$392/A1 U$$122/A2 U$$118/B1 U$$122/B2 VGND VGND VPWR VPWR U$$119/A sky130_fd_sc_hd__a22o_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater483 U$$3517/A2 VGND VGND VPWR VPWR U$$3549/A2 sky130_fd_sc_hd__buf_4
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_19_0 dadda_fa_7_19_0/A dadda_fa_7_19_0/B dadda_fa_7_19_0/CIN VGND VGND
+ VPWR VPWR _316_/D _187_/D sky130_fd_sc_hd__fa_1
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$129 U$$129/A U$$3/A VGND VGND VPWR VPWR U$$129/X sky130_fd_sc_hd__xor2_1
Xrepeater494 U$$3292/X VGND VGND VPWR VPWR U$$3378/A2 sky130_fd_sc_hd__buf_8
XU$$682_1840 VGND VGND VPWR VPWR U$$682_1840/HI U$$682/B1 sky130_fd_sc_hd__conb_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_426 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1007 input88/X VGND VGND VPWR VPWR U$$4452/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_110_0 dadda_fa_3_110_0/A U$$3286/X U$$3419/X VGND VGND VPWR VPWR dadda_fa_4_111_0/CIN
+ dadda_fa_4_110_1/CIN sky130_fd_sc_hd__fa_1
Xrepeater1018 U$$4450/A1 VGND VGND VPWR VPWR U$$1984/A1 sky130_fd_sc_hd__buf_6
Xrepeater1029 input85/X VGND VGND VPWR VPWR U$$3352/A1 sky130_fd_sc_hd__buf_8
XFILLER_181_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput220 c[67] VGND VGND VPWR VPWR input220/X sky130_fd_sc_hd__clkbuf_1
Xinput231 c[77] VGND VGND VPWR VPWR input231/X sky130_fd_sc_hd__buf_2
XFILLER_0_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput242 c[87] VGND VGND VPWR VPWR input242/X sky130_fd_sc_hd__clkbuf_2
Xdadda_fa_3_51_2 dadda_fa_3_51_2/A dadda_fa_3_51_2/B dadda_fa_3_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_1/A dadda_fa_4_51_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_0_67_2 U$$939/X U$$1072/X U$$1205/X VGND VGND VPWR VPWR dadda_fa_1_68_6/A
+ dadda_fa_1_67_8/A sky130_fd_sc_hd__fa_1
XFILLER_102_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_3_116_0_1874 VGND VGND VPWR VPWR dadda_ha_3_116_0/A dadda_ha_3_116_0_1874/LO
+ sky130_fd_sc_hd__conb_1
Xinput253 c[97] VGND VGND VPWR VPWR input253/X sky130_fd_sc_hd__clkbuf_4
XTAP_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_44_1 dadda_fa_3_44_1/A dadda_fa_3_44_1/B dadda_fa_3_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_0/CIN dadda_fa_4_44_2/A sky130_fd_sc_hd__fa_1
XTAP_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_21_0 dadda_fa_6_21_0/A dadda_fa_6_21_0/B dadda_fa_6_21_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_22_0/B dadda_fa_7_21_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_37_0 dadda_fa_3_37_0/A dadda_fa_3_37_0/B dadda_fa_3_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_0/B dadda_fa_4_37_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$780 final_adder.U$$780/A final_adder.U$$780/B VGND VGND VPWR VPWR
+ final_adder.U$$780/X sky130_fd_sc_hd__and2_1
XTAP_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$791 final_adder.U$$790/B final_adder.U$$711/X final_adder.U$$679/X
+ VGND VGND VPWR VPWR final_adder.U$$791/X sky130_fd_sc_hd__a21o_1
XU$$630 U$$630/A1 U$$672/A2 U$$630/B1 U$$668/B2 VGND VGND VPWR VPWR U$$631/A sky130_fd_sc_hd__a22o_1
XFILLER_84_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$641 U$$641/A U$$651/B VGND VGND VPWR VPWR U$$641/X sky130_fd_sc_hd__xor2_1
XU$$652 U$$652/A1 U$$652/A2 U$$654/A1 U$$652/B2 VGND VGND VPWR VPWR U$$653/A sky130_fd_sc_hd__a22o_1
XU$$663 U$$663/A U$$673/B VGND VGND VPWR VPWR U$$663/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$674 U$$674/A1 U$$678/A2 U$$676/A1 U$$553/X VGND VGND VPWR VPWR U$$675/A sky130_fd_sc_hd__a22o_1
XU$$685 U$$685/A VGND VGND VPWR VPWR U$$685/Y sky130_fd_sc_hd__inv_1
XU$$696 U$$696/A U$$784/B VGND VGND VPWR VPWR U$$696/X sky130_fd_sc_hd__xor2_1
XFILLER_16_275 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_971 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_96_4 U$$4056/X U$$4189/X U$$4322/X VGND VGND VPWR VPWR dadda_fa_3_97_1/CIN
+ dadda_fa_3_96_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1530 U$$43/B VGND VGND VPWR VPWR U$$9/B sky130_fd_sc_hd__buf_4
Xrepeater1541 U$$3960/B1 VGND VGND VPWR VPWR U$$4236/A1 sky130_fd_sc_hd__buf_6
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1552 U$$3960/A1 VGND VGND VPWR VPWR U$$4508/A1 sky130_fd_sc_hd__buf_8
Xrepeater1563 U$$118/B1 VGND VGND VPWR VPWR U$$942/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_89_3 input244/X dadda_fa_2_89_3/B dadda_fa_2_89_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_90_1/B dadda_fa_3_89_3/B sky130_fd_sc_hd__fa_2
XFILLER_126_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1574 U$$2445/B1 VGND VGND VPWR VPWR U$$940/A1 sky130_fd_sc_hd__buf_4
XFILLER_67_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1585 U$$4361/B1 VGND VGND VPWR VPWR U$$4500/A1 sky130_fd_sc_hd__buf_6
XFILLER_67_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1596 input112/X VGND VGND VPWR VPWR U$$3946/B1 sky130_fd_sc_hd__buf_4
XFILLER_141_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4417_1785 VGND VGND VPWR VPWR U$$4417_1785/HI U$$4417/B sky130_fd_sc_hd__conb_1
Xdadda_fa_5_59_1 dadda_fa_5_59_1/A dadda_fa_5_59_1/B dadda_fa_5_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_60_0/B dadda_fa_7_59_0/A sky130_fd_sc_hd__fa_1
XFILLER_58_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_105_1 U$$3276/X U$$3409/X U$$3542/X VGND VGND VPWR VPWR dadda_fa_3_106_3/B
+ dadda_fa_4_105_0/A sky130_fd_sc_hd__fa_1
XFILLER_39_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2070 U$$2070/A U$$2100/B VGND VGND VPWR VPWR U$$2070/X sky130_fd_sc_hd__xor2_1
XU$$2081 U$$2492/A1 U$$2091/A2 U$$2220/A1 U$$2091/B2 VGND VGND VPWR VPWR U$$2082/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2092 U$$2092/A U$$2092/B VGND VGND VPWR VPWR U$$2092/X sky130_fd_sc_hd__xor2_1
XFILLER_165_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1380 U$$2202/A1 U$$1404/A2 U$$2202/B1 U$$1404/B2 VGND VGND VPWR VPWR U$$1381/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1391 U$$1391/A U$$1399/B VGND VGND VPWR VPWR U$$1391/X sky130_fd_sc_hd__xor2_1
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_478 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_84_2 U$$2170/X U$$2303/X U$$2436/X VGND VGND VPWR VPWR dadda_fa_2_85_2/CIN
+ dadda_fa_2_84_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_61_1 dadda_fa_4_61_1/A dadda_fa_4_61_1/B dadda_fa_4_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/B dadda_fa_5_61_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_77_1 U$$1757/X U$$1890/X U$$2023/X VGND VGND VPWR VPWR dadda_fa_2_78_0/CIN
+ dadda_fa_2_77_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_54_0 dadda_fa_4_54_0/A dadda_fa_4_54_0/B dadda_fa_4_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/A dadda_fa_5_54_1/A sky130_fd_sc_hd__fa_1
XTAP_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1018 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_372_ _373_/CLK _372_/D VGND VGND VPWR VPWR _372_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_99_2 dadda_fa_3_99_2/A dadda_fa_3_99_2/B dadda_fa_3_99_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_1/A dadda_fa_4_99_2/B sky130_fd_sc_hd__fa_1
XFILLER_6_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_69_0 dadda_fa_6_69_0/A dadda_fa_6_69_0/B dadda_fa_6_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_70_0/B dadda_fa_7_69_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_205_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_72_0 dadda_fa_0_72_0/A U$$683/X U$$816/X VGND VGND VPWR VPWR dadda_fa_1_73_7/A
+ dadda_fa_1_72_8/A sky130_fd_sc_hd__fa_1
XFILLER_95_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$460 U$$460/A U$$492/B VGND VGND VPWR VPWR U$$460/X sky130_fd_sc_hd__xor2_1
XU$$471 U$$745/A1 U$$473/A2 U$$882/B1 U$$473/B2 VGND VGND VPWR VPWR U$$472/A sky130_fd_sc_hd__a22o_1
XFILLER_44_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$482 U$$482/A U$$484/B VGND VGND VPWR VPWR U$$482/X sky130_fd_sc_hd__xor2_1
XU$$493 U$$630/A1 U$$537/A2 U$$630/B1 U$$537/B2 VGND VGND VPWR VPWR U$$494/A sky130_fd_sc_hd__a22o_1
XFILLER_204_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_271 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_94_1 U$$3121/X U$$3254/X U$$3387/X VGND VGND VPWR VPWR dadda_fa_3_95_0/CIN
+ dadda_fa_3_94_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_71_0 dadda_fa_5_71_0/A dadda_fa_5_71_0/B dadda_fa_5_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_72_0/A dadda_fa_6_71_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_87_0 U$$3639/X U$$3772/X U$$3905/X VGND VGND VPWR VPWR dadda_fa_3_88_0/B
+ dadda_fa_3_87_2/B sky130_fd_sc_hd__fa_1
Xrepeater1360 U$$2716/B VGND VGND VPWR VPWR U$$2658/B sky130_fd_sc_hd__buf_6
XFILLER_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1371 U$$2569/B VGND VGND VPWR VPWR U$$2543/B sky130_fd_sc_hd__buf_8
XFILLER_114_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1382 U$$808/B VGND VGND VPWR VPWR U$$796/B sky130_fd_sc_hd__buf_6
Xrepeater1393 U$$2253/B VGND VGND VPWR VPWR U$$2227/B sky130_fd_sc_hd__buf_8
XFILLER_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_70_8 dadda_fa_1_70_8/A dadda_fa_1_70_8/B dadda_fa_1_70_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_71_3/A dadda_fa_3_70_0/A sky130_fd_sc_hd__fa_1
XFILLER_114_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_63_7 dadda_fa_1_63_7/A dadda_fa_1_63_7/B dadda_fa_1_63_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_2/CIN dadda_fa_2_63_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_56_6 U$$3577/X U$$3710/X U$$3843/X VGND VGND VPWR VPWR dadda_fa_2_57_2/B
+ dadda_fa_2_56_5/B sky130_fd_sc_hd__fa_1
XFILLER_28_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_49_5 U$$2100/X U$$2233/X U$$2366/X VGND VGND VPWR VPWR dadda_fa_2_50_2/B
+ dadda_fa_2_49_5/B sky130_fd_sc_hd__fa_1
XFILLER_82_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_8_0 dadda_fa_7_8_0/A dadda_fa_7_8_0/B dadda_fa_7_8_0/CIN VGND VGND VPWR
+ VPWR _305_/D _176_/D sky130_fd_sc_hd__fa_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_532 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_86_0 dadda_fa_7_86_0/A dadda_fa_7_86_0/B dadda_fa_7_86_0/CIN VGND VGND
+ VPWR VPWR _383_/D _254_/D sky130_fd_sc_hd__fa_1
XFILLER_148_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4208 U$$4343/B1 U$$4210/A2 U$$4210/A1 U$$4210/B2 VGND VGND VPWR VPWR U$$4209/A
+ sky130_fd_sc_hd__a22o_1
XU$$4219 U$$4219/A U$$4247/A VGND VGND VPWR VPWR U$$4219/X sky130_fd_sc_hd__xor2_1
XU$$3507 U$$3644/A1 U$$3429/X U$$3644/B1 U$$3430/X VGND VGND VPWR VPWR U$$3508/A sky130_fd_sc_hd__a22o_1
XFILLER_74_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3518 U$$3518/A U$$3518/B VGND VGND VPWR VPWR U$$3518/X sky130_fd_sc_hd__xor2_1
XFILLER_100_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_101_0 dadda_fa_6_101_0/A dadda_fa_6_101_0/B dadda_fa_6_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_102_0/B dadda_fa_7_101_0/CIN sky130_fd_sc_hd__fa_1
XU$$3529 U$$3801/B1 U$$3549/A2 U$$4077/B1 U$$3549/B2 VGND VGND VPWR VPWR U$$3530/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2806 U$$3078/B1 U$$2810/A2 U$$3902/B1 U$$2810/B2 VGND VGND VPWR VPWR U$$2807/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_100 _346_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2817 U$$2817/A U$$2817/B VGND VGND VPWR VPWR U$$2817/X sky130_fd_sc_hd__xor2_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2828 U$$3648/B1 U$$2828/A2 U$$3378/A1 U$$2828/B2 VGND VGND VPWR VPWR U$$2829/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2839 U$$2839/A U$$2845/B VGND VGND VPWR VPWR U$$2839/X sky130_fd_sc_hd__xor2_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_122 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 U$$3356/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_144 U$$1746/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 U$$2737/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_177 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_188 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_199 _199_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_355_ _355_/CLK _355_/D VGND VGND VPWR VPWR _355_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_286_ _417_/CLK _286_/D VGND VGND VPWR VPWR _286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_66_5 dadda_fa_2_66_5/A dadda_fa_2_66_5/B dadda_fa_2_66_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_67_2/A dadda_fa_4_66_0/A sky130_fd_sc_hd__fa_2
XFILLER_111_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_59_4 dadda_fa_2_59_4/A dadda_fa_2_59_4/B dadda_fa_2_59_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_1/CIN dadda_fa_3_59_3/CIN sky130_fd_sc_hd__fa_1
XTAP_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 a[14] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$290 U$$16/A1 U$$302/A2 U$$703/A1 U$$302/B2 VGND VGND VPWR VPWR U$$291/A sky130_fd_sc_hd__a22o_1
XFILLER_36_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$4 _300_/Q _172_/Q VGND VGND VPWR VPWR final_adder.U$$4/COUT final_adder.U$$4/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_69_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput310 output310/A VGND VGND VPWR VPWR o[32] sky130_fd_sc_hd__buf_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput321 output321/A VGND VGND VPWR VPWR o[42] sky130_fd_sc_hd__buf_2
Xoutput332 output332/A VGND VGND VPWR VPWR o[52] sky130_fd_sc_hd__buf_2
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 output343/A VGND VGND VPWR VPWR o[62] sky130_fd_sc_hd__buf_2
XFILLER_114_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput354 output354/A VGND VGND VPWR VPWR o[72] sky130_fd_sc_hd__buf_2
Xoutput365 output365/A VGND VGND VPWR VPWR o[82] sky130_fd_sc_hd__buf_2
Xoutput376 output376/A VGND VGND VPWR VPWR o[92] sky130_fd_sc_hd__buf_2
Xrepeater1190 U$$711/B1 VGND VGND VPWR VPWR U$$850/A1 sky130_fd_sc_hd__buf_6
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_61_4 U$$3587/X U$$3720/X U$$3853/X VGND VGND VPWR VPWR dadda_fa_2_62_1/CIN
+ dadda_fa_2_61_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_45_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_3 U$$1977/X U$$2110/X U$$2243/X VGND VGND VPWR VPWR dadda_fa_2_55_1/B
+ dadda_fa_2_54_4/B sky130_fd_sc_hd__fa_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_31_2 dadda_fa_4_31_2/A dadda_fa_4_31_2/B dadda_fa_4_31_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_32_0/CIN dadda_fa_5_31_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_47_2 U$$899/X U$$1032/X U$$1165/X VGND VGND VPWR VPWR dadda_fa_2_48_2/A
+ dadda_fa_2_47_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_56_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_24_1 dadda_fa_4_24_1/A dadda_fa_4_24_1/B dadda_fa_4_24_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/B dadda_fa_5_24_1/B sky130_fd_sc_hd__fa_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_17_0 U$$706/X U$$839/X U$$972/X VGND VGND VPWR VPWR dadda_fa_5_18_0/A
+ dadda_fa_5_17_1/A sky130_fd_sc_hd__fa_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_868 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_69_3 dadda_fa_3_69_3/A dadda_fa_3_69_3/B dadda_fa_3_69_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_70_1/B dadda_fa_4_69_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4005 U$$4005/A1 U$$4011/A2 U$$4005/B1 U$$4011/B2 VGND VGND VPWR VPWR U$$4006/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4016 U$$4016/A U$$4080/B VGND VGND VPWR VPWR U$$4016/X sky130_fd_sc_hd__xor2_1
XFILLER_76_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4027 U$$4027/A1 U$$4043/A2 U$$4029/A1 U$$4043/B2 VGND VGND VPWR VPWR U$$4028/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4038 U$$4038/A U$$4109/A VGND VGND VPWR VPWR U$$4038/X sky130_fd_sc_hd__xor2_1
XU$$3304 U$$3578/A1 U$$3394/A2 U$$3578/B1 U$$3394/B2 VGND VGND VPWR VPWR U$$3305/A
+ sky130_fd_sc_hd__a22o_1
XU$$4049 input92/X U$$4079/A2 U$$4049/B1 U$$4079/B2 VGND VGND VPWR VPWR U$$4050/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3315 U$$3315/A U$$3321/B VGND VGND VPWR VPWR U$$3315/X sky130_fd_sc_hd__xor2_1
XU$$3326 U$$3737/A1 U$$3348/A2 U$$3737/B1 U$$3346/B2 VGND VGND VPWR VPWR U$$3327/A
+ sky130_fd_sc_hd__a22o_1
XU$$3337 U$$3337/A U$$3377/B VGND VGND VPWR VPWR U$$3337/X sky130_fd_sc_hd__xor2_1
XFILLER_47_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2603 U$$2603/A VGND VGND VPWR VPWR U$$2603/Y sky130_fd_sc_hd__inv_1
XFILLER_202_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3348 U$$3483/B1 U$$3348/A2 U$$3348/B1 U$$3394/B2 VGND VGND VPWR VPWR U$$3349/A
+ sky130_fd_sc_hd__a22o_1
XU$$2614 U$$2614/A U$$2624/B VGND VGND VPWR VPWR U$$2614/X sky130_fd_sc_hd__xor2_1
XU$$3359 U$$3359/A U$$3425/A VGND VGND VPWR VPWR U$$3359/X sky130_fd_sc_hd__xor2_1
XU$$2625 U$$2625/A1 U$$2625/A2 U$$2625/B1 U$$2625/B2 VGND VGND VPWR VPWR U$$2626/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2636 U$$2636/A U$$2650/B VGND VGND VPWR VPWR U$$2636/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2647 U$$4015/B1 U$$2727/A2 U$$4019/A1 U$$2727/B2 VGND VGND VPWR VPWR U$$2648/A
+ sky130_fd_sc_hd__a22o_1
XU$$1902 U$$1902/A U$$1914/B VGND VGND VPWR VPWR U$$1902/X sky130_fd_sc_hd__xor2_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2658 U$$2658/A U$$2658/B VGND VGND VPWR VPWR U$$2658/X sky130_fd_sc_hd__xor2_1
XU$$1913 U$$4516/A1 U$$1913/A2 U$$4516/B1 U$$1786/X VGND VGND VPWR VPWR U$$1914/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1924 U$$1924/A1 U$$1960/A2 U$$2198/B1 U$$1960/B2 VGND VGND VPWR VPWR U$$1925/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2669 U$$3078/B1 U$$2691/A2 U$$3356/A1 U$$2691/B2 VGND VGND VPWR VPWR U$$2670/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1935 U$$1935/A U$$1971/B VGND VGND VPWR VPWR U$$1935/X sky130_fd_sc_hd__xor2_1
XU$$1946 U$$2220/A1 U$$1960/A2 U$$3727/B1 U$$1960/B2 VGND VGND VPWR VPWR U$$1947/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1957 U$$1957/A U$$1993/B VGND VGND VPWR VPWR U$$1957/X sky130_fd_sc_hd__xor2_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1968 U$$50/A1 U$$1970/A2 U$$3749/B1 U$$1970/B2 VGND VGND VPWR VPWR U$$1969/A sky130_fd_sc_hd__a22o_1
X_407_ _407_/CLK _407_/D VGND VGND VPWR VPWR _407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1979 U$$1979/A U$$2017/B VGND VGND VPWR VPWR U$$1979/X sky130_fd_sc_hd__xor2_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_986 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_338_ _351_/CLK _338_/D VGND VGND VPWR VPWR _338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_269_ _397_/CLK _269_/D VGND VGND VPWR VPWR _269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_426 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_278 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_71_3 dadda_fa_2_71_3/A dadda_fa_2_71_3/B dadda_fa_2_71_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/B dadda_fa_3_71_3/B sky130_fd_sc_hd__fa_1
XFILLER_124_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_64_2 dadda_fa_2_64_2/A dadda_fa_2_64_2/B dadda_fa_2_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/A dadda_fa_3_64_3/A sky130_fd_sc_hd__fa_1
Xrepeater802 U$$2449/B2 VGND VGND VPWR VPWR U$$2435/B2 sky130_fd_sc_hd__buf_6
XFILLER_110_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$609 final_adder.U$$608/B final_adder.U$$493/X final_adder.U$$485/X
+ VGND VGND VPWR VPWR final_adder.U$$609/X sky130_fd_sc_hd__a21o_1
Xrepeater813 U$$2197/X VGND VGND VPWR VPWR U$$2302/B2 sky130_fd_sc_hd__buf_6
XFILLER_96_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_41_1 dadda_fa_5_41_1/A dadda_fa_5_41_1/B dadda_fa_5_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_42_0/B dadda_fa_7_41_0/A sky130_fd_sc_hd__fa_2
Xrepeater824 U$$2016/B2 VGND VGND VPWR VPWR U$$1990/B2 sky130_fd_sc_hd__buf_8
XFILLER_110_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_57_1 dadda_fa_2_57_1/A dadda_fa_2_57_1/B dadda_fa_2_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_0/CIN dadda_fa_3_57_2/CIN sky130_fd_sc_hd__fa_2
Xrepeater835 U$$1903/B2 VGND VGND VPWR VPWR U$$1915/B2 sky130_fd_sc_hd__buf_8
Xrepeater846 U$$1649/X VGND VGND VPWR VPWR U$$1770/B2 sky130_fd_sc_hd__buf_6
XFILLER_42_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater857 U$$209/B2 VGND VGND VPWR VPWR U$$175/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_34_0 dadda_fa_5_34_0/A dadda_fa_5_34_0/B dadda_fa_5_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_35_0/A dadda_fa_6_34_0/CIN sky130_fd_sc_hd__fa_1
XU$$20 U$$20/A1 U$$42/A2 U$$22/A1 U$$42/B2 VGND VGND VPWR VPWR U$$21/A sky130_fd_sc_hd__a22o_1
Xrepeater868 U$$1470/B2 VGND VGND VPWR VPWR U$$1462/B2 sky130_fd_sc_hd__buf_4
XFILLER_110_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater879 U$$1190/B2 VGND VGND VPWR VPWR U$$1136/B2 sky130_fd_sc_hd__buf_4
XU$$31 U$$31/A U$$51/B VGND VGND VPWR VPWR U$$31/X sky130_fd_sc_hd__xor2_1
XFILLER_53_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$42 U$$42/A1 U$$42/A2 U$$44/A1 U$$42/B2 VGND VGND VPWR VPWR U$$43/A sky130_fd_sc_hd__a22o_1
XU$$53 U$$53/A U$$81/B VGND VGND VPWR VPWR U$$53/X sky130_fd_sc_hd__xor2_1
XU$$64 U$$64/A1 U$$98/A2 U$$66/A1 U$$98/B2 VGND VGND VPWR VPWR U$$65/A sky130_fd_sc_hd__a22o_1
XFILLER_65_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3860 U$$4269/B1 U$$3874/A2 U$$4408/B1 U$$3874/B2 VGND VGND VPWR VPWR U$$3861/A
+ sky130_fd_sc_hd__a22o_1
XU$$75 U$$75/A U$$81/B VGND VGND VPWR VPWR U$$75/X sky130_fd_sc_hd__xor2_1
XU$$3871 U$$3871/A U$$3903/B VGND VGND VPWR VPWR U$$3871/X sky130_fd_sc_hd__xor2_1
XFILLER_53_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3882 U$$4019/A1 U$$3926/A2 U$$3882/B1 U$$3926/B2 VGND VGND VPWR VPWR U$$3883/A
+ sky130_fd_sc_hd__a22o_1
XU$$86 U$$86/A1 U$$94/A2 U$$88/A1 U$$94/B2 VGND VGND VPWR VPWR U$$87/A sky130_fd_sc_hd__a22o_1
XU$$97 U$$97/A U$$99/B VGND VGND VPWR VPWR U$$97/X sky130_fd_sc_hd__xor2_1
XFILLER_64_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3893 U$$3893/A U$$3909/B VGND VGND VPWR VPWR U$$3893/X sky130_fd_sc_hd__xor2_1
XFILLER_52_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_11 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _336_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_33 _339_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_44 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_55 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_66 _342_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_398 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_99 _346_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_79_2 dadda_fa_4_79_2/A dadda_fa_4_79_2/B dadda_fa_4_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_80_0/CIN dadda_fa_5_79_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_173_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_941 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_49_0 dadda_fa_7_49_0/A dadda_fa_7_49_0/B dadda_fa_7_49_0/CIN VGND VGND
+ VPWR VPWR _346_/D _217_/D sky130_fd_sc_hd__fa_2
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1039 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_52_0 U$$377/X U$$510/X U$$643/X VGND VGND VPWR VPWR dadda_fa_2_53_0/B
+ dadda_fa_2_52_3/B sky130_fd_sc_hd__fa_1
XFILLER_28_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1209 U$$1209/A U$$1209/B VGND VGND VPWR VPWR U$$1209/X sky130_fd_sc_hd__xor2_1
XFILLER_203_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$1003 final_adder.U$$232/A final_adder.U$$733/X final_adder.U$$233/A2
+ VGND VGND VPWR VPWR final_adder.U$$1047/B sky130_fd_sc_hd__a21o_1
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1025 final_adder.U$$1/SUM final_adder.U$$255/A2 VGND VGND VPWR VPWR
+ output296/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1036 final_adder.U$$242/A final_adder.U$$623/X VGND VGND VPWR VPWR
+ output288/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1047 final_adder.U$$232/B final_adder.U$$1047/B VGND VGND VPWR VPWR
+ output300/A sky130_fd_sc_hd__xor2_1
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1058 final_adder.U$$220/A final_adder.U$$833/X VGND VGND VPWR VPWR
+ output312/A sky130_fd_sc_hd__xor2_1
XFILLER_165_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1069 final_adder.U$$210/B final_adder.U$$981/X VGND VGND VPWR VPWR
+ output324/A sky130_fd_sc_hd__xor2_1
XFILLER_164_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_81_2 dadda_fa_3_81_2/A dadda_fa_3_81_2/B dadda_fa_3_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_1/A dadda_fa_4_81_2/B sky130_fd_sc_hd__fa_1
XFILLER_112_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_74_1 dadda_fa_3_74_1/A dadda_fa_3_74_1/B dadda_fa_3_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_0/CIN dadda_fa_4_74_2/A sky130_fd_sc_hd__fa_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_51_0 dadda_fa_6_51_0/A dadda_fa_6_51_0/B dadda_fa_6_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_52_0/B dadda_fa_7_51_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_26_1226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_67_0 dadda_fa_3_67_0/A dadda_fa_3_67_0/B dadda_fa_3_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_0/B dadda_fa_4_67_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3101 U$$3101/A U$$3109/B VGND VGND VPWR VPWR U$$3101/X sky130_fd_sc_hd__xor2_1
XFILLER_94_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3112 U$$3112/A1 U$$3018/X U$$3114/A1 U$$3019/X VGND VGND VPWR VPWR U$$3113/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_110_2 dadda_fa_4_110_2/A dadda_fa_4_110_2/B dadda_ha_3_110_3/SUM VGND
+ VGND VPWR VPWR dadda_fa_5_111_0/CIN dadda_fa_5_110_1/CIN sky130_fd_sc_hd__fa_1
XU$$3123 U$$3123/A U$$3133/B VGND VGND VPWR VPWR U$$3123/X sky130_fd_sc_hd__xor2_1
XU$$3134 U$$3545/A1 U$$3148/A2 U$$3684/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3135/A
+ sky130_fd_sc_hd__a22o_1
XU$$3145 U$$3145/A U$$3150/A VGND VGND VPWR VPWR U$$3145/X sky130_fd_sc_hd__xor2_1
XU$$2400 U$$2400/A U$$2442/B VGND VGND VPWR VPWR U$$2400/X sky130_fd_sc_hd__xor2_1
XFILLER_47_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2411 U$$3368/B1 U$$2435/A2 U$$3646/A1 U$$2435/B2 VGND VGND VPWR VPWR U$$2412/A
+ sky130_fd_sc_hd__a22o_1
XU$$3156 U$$3154/B U$$3151/A input41/X U$$3151/Y VGND VGND VPWR VPWR U$$3156/X sky130_fd_sc_hd__a22o_4
XFILLER_98_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_103_1 dadda_fa_4_103_1/A dadda_fa_4_103_1/B dadda_fa_4_103_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/B dadda_fa_5_103_1/B sky130_fd_sc_hd__fa_1
XU$$2422 U$$2422/A U$$2454/B VGND VGND VPWR VPWR U$$2422/X sky130_fd_sc_hd__xor2_1
XFILLER_207_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3167 input109/X U$$3187/A2 U$$3578/B1 U$$3187/B2 VGND VGND VPWR VPWR U$$3168/A
+ sky130_fd_sc_hd__a22o_1
XU$$3178 U$$3178/A U$$3264/B VGND VGND VPWR VPWR U$$3178/X sky130_fd_sc_hd__xor2_1
XU$$2433 U$$3116/B1 U$$2449/A2 U$$2981/B1 U$$2449/B2 VGND VGND VPWR VPWR U$$2434/A
+ sky130_fd_sc_hd__a22o_1
XU$$2444 U$$2444/A U$$2466/A VGND VGND VPWR VPWR U$$2444/X sky130_fd_sc_hd__xor2_1
XU$$3189 U$$860/A1 U$$3207/A2 U$$3737/B1 U$$3207/B2 VGND VGND VPWR VPWR U$$3190/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2455 U$$3960/B1 U$$2459/A2 U$$3416/A1 U$$2459/B2 VGND VGND VPWR VPWR U$$2456/A
+ sky130_fd_sc_hd__a22o_1
XU$$1710 U$$1984/A1 U$$1750/A2 U$$342/A1 U$$1750/B2 VGND VGND VPWR VPWR U$$1711/A
+ sky130_fd_sc_hd__a22o_1
XU$$2466 U$$2466/A VGND VGND VPWR VPWR U$$2466/Y sky130_fd_sc_hd__inv_1
XU$$1721 U$$1721/A U$$1721/B VGND VGND VPWR VPWR U$$1721/X sky130_fd_sc_hd__xor2_1
XU$$1732 U$$3376/A1 U$$1736/A2 U$$3102/B1 U$$1736/B2 VGND VGND VPWR VPWR U$$1733/A
+ sky130_fd_sc_hd__a22o_1
XU$$2477 U$$2477/A U$$2525/B VGND VGND VPWR VPWR U$$2477/X sky130_fd_sc_hd__xor2_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1743 U$$1743/A U$$1780/A VGND VGND VPWR VPWR U$$1743/X sky130_fd_sc_hd__xor2_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2488 U$$2625/A1 U$$2490/A2 U$$2625/B1 U$$2490/B2 VGND VGND VPWR VPWR U$$2489/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2499 U$$2499/A U$$2543/B VGND VGND VPWR VPWR U$$2499/X sky130_fd_sc_hd__xor2_1
XU$$1754 U$$384/A1 U$$1764/A2 U$$521/B1 U$$1764/B2 VGND VGND VPWR VPWR U$$1755/A sky130_fd_sc_hd__a22o_1
XU$$1765 U$$1765/A U$$1765/B VGND VGND VPWR VPWR U$$1765/X sky130_fd_sc_hd__xor2_1
XFILLER_203_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1776 U$$4516/A1 U$$1648/X U$$4516/B1 U$$1649/X VGND VGND VPWR VPWR U$$1777/A sky130_fd_sc_hd__a22o_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1787 U$$1787/A1 U$$1819/A2 U$$2198/B1 U$$1819/B2 VGND VGND VPWR VPWR U$$1788/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1798 U$$1798/A U$$1832/B VGND VGND VPWR VPWR U$$1798/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_124_0 dadda_fa_7_124_0/A dadda_fa_7_124_0/B dadda_fa_7_124_0/CIN VGND
+ VGND VPWR VPWR _421_/D _292_/D sky130_fd_sc_hd__fa_2
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_clk _385_/CLK VGND VGND VPWR VPWR _421_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_147_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput20 a[27] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__buf_4
Xinput31 a[37] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__buf_4
XFILLER_190_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput42 a[47] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 a[57] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput64 a[9] VGND VGND VPWR VPWR U$$683/B sky130_fd_sc_hd__buf_6
Xinput75 b[19] VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__buf_12
Xdadda_fa_5_89_1 dadda_fa_5_89_1/A dadda_fa_5_89_1/B dadda_fa_5_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_90_0/B dadda_fa_7_89_0/A sky130_fd_sc_hd__fa_1
Xinput86 b[29] VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__buf_6
XFILLER_115_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput97 b[39] VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__buf_6
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$406 final_adder.U$$410/B final_adder.U$$406/B VGND VGND VPWR VPWR
+ final_adder.U$$530/B sky130_fd_sc_hd__and2_1
Xrepeater610 U$$209/A2 VGND VGND VPWR VPWR U$$175/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_97_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$417 final_adder.U$$416/B final_adder.U$$295/X final_adder.U$$291/X
+ VGND VGND VPWR VPWR final_adder.U$$417/X sky130_fd_sc_hd__a21o_1
Xrepeater621 U$$1470/A2 VGND VGND VPWR VPWR U$$1462/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$428 final_adder.U$$432/B final_adder.U$$428/B VGND VGND VPWR VPWR
+ final_adder.U$$552/B sky130_fd_sc_hd__and2_1
XFILLER_96_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater632 U$$1190/A2 VGND VGND VPWR VPWR U$$1136/A2 sky130_fd_sc_hd__buf_4
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$439 final_adder.U$$438/B final_adder.U$$317/X final_adder.U$$313/X
+ VGND VGND VPWR VPWR final_adder.U$$439/X sky130_fd_sc_hd__a21o_1
XFILLER_38_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater643 U$$1057/B2 VGND VGND VPWR VPWR U$$997/B2 sky130_fd_sc_hd__buf_4
Xrepeater654 U$$827/X VGND VGND VPWR VPWR U$$938/B2 sky130_fd_sc_hd__buf_4
XFILLER_42_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater665 U$$652/B2 VGND VGND VPWR VPWR U$$578/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_72_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater676 U$$4373/B2 VGND VGND VPWR VPWR U$$4369/B2 sky130_fd_sc_hd__buf_4
Xrepeater687 U$$4176/B2 VGND VGND VPWR VPWR U$$4164/B2 sky130_fd_sc_hd__buf_4
XFILLER_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4380 U$$4380/A U$$4382/B VGND VGND VPWR VPWR U$$4380/X sky130_fd_sc_hd__xor2_1
Xrepeater698 U$$4107/B2 VGND VGND VPWR VPWR U$$4103/B2 sky130_fd_sc_hd__buf_4
XU$$4391 U$$4391/A U$$4391/B VGND VGND VPWR VPWR U$$4391/X sky130_fd_sc_hd__xor2_1
XFILLER_25_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3690 U$$4099/B1 U$$3696/A2 U$$4240/A1 U$$3696/B2 VGND VGND VPWR VPWR U$$3691/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_clk _255_/CLK VGND VGND VPWR VPWR _417_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_91_1 dadda_fa_4_91_1/A dadda_fa_4_91_1/B dadda_fa_4_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_92_0/B dadda_fa_5_91_1/B sky130_fd_sc_hd__fa_1
XFILLER_181_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_84_0 dadda_fa_4_84_0/A dadda_fa_4_84_0/B dadda_fa_4_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/A dadda_fa_5_84_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_105_3 dadda_fa_3_105_3/A dadda_fa_3_105_3/B dadda_fa_3_105_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_106_1/B dadda_fa_4_105_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_101_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$951 final_adder.U$$180/A final_adder.U$$889/X final_adder.U$$951/B1
+ VGND VGND VPWR VPWR final_adder.U$$951/X sky130_fd_sc_hd__a21o_1
XTAP_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$801 U$$938/A1 U$$805/A2 U$$940/A1 U$$805/B2 VGND VGND VPWR VPWR U$$802/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$973 final_adder.U$$202/A final_adder.U$$815/X final_adder.U$$973/B1
+ VGND VGND VPWR VPWR final_adder.U$$973/X sky130_fd_sc_hd__a21o_1
XU$$812 U$$812/A U$$821/A VGND VGND VPWR VPWR U$$812/X sky130_fd_sc_hd__xor2_1
XTAP_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$823 input4/X VGND VGND VPWR VPWR U$$825/B sky130_fd_sc_hd__inv_1
XFILLER_95_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$995 final_adder.U$$224/A final_adder.U$$725/X final_adder.U$$995/B1
+ VGND VGND VPWR VPWR final_adder.U$$995/X sky130_fd_sc_hd__a21o_1
XU$$834 U$$969/B1 U$$906/A2 U$$836/A1 U$$906/B2 VGND VGND VPWR VPWR U$$835/A sky130_fd_sc_hd__a22o_1
XFILLER_17_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$845 U$$845/A U$$847/B VGND VGND VPWR VPWR U$$845/X sky130_fd_sc_hd__xor2_1
XFILLER_21_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$856 U$$993/A1 U$$892/A2 U$$993/B1 U$$892/B2 VGND VGND VPWR VPWR U$$857/A sky130_fd_sc_hd__a22o_1
XFILLER_189_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_969 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$867 U$$867/A U$$877/B VGND VGND VPWR VPWR U$$867/X sky130_fd_sc_hd__xor2_1
XU$$1006 U$$1006/A U$$996/B VGND VGND VPWR VPWR U$$1006/X sky130_fd_sc_hd__xor2_1
XU$$1017 U$$58/A1 U$$993/A2 U$$60/A1 U$$993/B2 VGND VGND VPWR VPWR U$$1018/A sky130_fd_sc_hd__a22o_1
XU$$878 U$$56/A1 U$$882/A2 U$$878/B1 U$$882/B2 VGND VGND VPWR VPWR U$$879/A sky130_fd_sc_hd__a22o_1
XU$$1028 U$$1028/A U$$1076/B VGND VGND VPWR VPWR U$$1028/X sky130_fd_sc_hd__xor2_1
XU$$889 U$$889/A U$$929/B VGND VGND VPWR VPWR U$$889/X sky130_fd_sc_hd__xor2_1
XU$$1039 U$$902/A1 U$$979/A2 U$$82/A1 U$$979/B2 VGND VGND VPWR VPWR U$$1040/A sky130_fd_sc_hd__a22o_1
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_clk _380_/CLK VGND VGND VPWR VPWR _401_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_6_99_0 dadda_fa_6_99_0/A dadda_fa_6_99_0/B dadda_fa_6_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_100_0/B dadda_fa_7_99_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_157_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1701 U$$912/A1 VGND VGND VPWR VPWR U$$773/B1 sky130_fd_sc_hd__buf_6
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1048 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_41_4 dadda_fa_2_41_4/A dadda_fa_2_41_4/B dadda_fa_2_41_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_42_1/CIN dadda_fa_3_41_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_34_3 U$$1538/X U$$1671/X U$$1804/X VGND VGND VPWR VPWR dadda_fa_3_35_1/B
+ dadda_fa_3_34_3/B sky130_fd_sc_hd__fa_1
XFILLER_208_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2230 U$$4011/A1 U$$2252/A2 U$$4011/B1 U$$2252/B2 VGND VGND VPWR VPWR U$$2231/A
+ sky130_fd_sc_hd__a22o_1
XU$$2241 U$$2241/A U$$2285/B VGND VGND VPWR VPWR U$$2241/X sky130_fd_sc_hd__xor2_1
XFILLER_207_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2252 U$$3483/B1 U$$2252/A2 U$$610/A1 U$$2252/B2 VGND VGND VPWR VPWR U$$2253/A
+ sky130_fd_sc_hd__a22o_1
XU$$2263 U$$2263/A U$$2309/B VGND VGND VPWR VPWR U$$2263/X sky130_fd_sc_hd__xor2_1
XU$$2274 U$$3368/B1 U$$2302/A2 U$$3646/A1 U$$2302/B2 VGND VGND VPWR VPWR U$$2275/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1540 U$$1540/A U$$1574/B VGND VGND VPWR VPWR U$$1540/X sky130_fd_sc_hd__xor2_1
XU$$2285 U$$2285/A U$$2285/B VGND VGND VPWR VPWR U$$2285/X sky130_fd_sc_hd__xor2_1
XU$$1551 U$$727/B1 U$$1557/A2 U$$594/A1 U$$1557/B2 VGND VGND VPWR VPWR U$$1552/A sky130_fd_sc_hd__a22o_1
XU$$2296 U$$3116/B1 U$$2316/A2 U$$2981/B1 U$$2316/B2 VGND VGND VPWR VPWR U$$2297/A
+ sky130_fd_sc_hd__a22o_1
XU$$1562 U$$1562/A U$$1592/B VGND VGND VPWR VPWR U$$1562/X sky130_fd_sc_hd__xor2_1
XFILLER_22_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1573 U$$1984/A1 U$$1575/A2 U$$342/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1574/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_clk _227_/CLK VGND VGND VPWR VPWR _355_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1584 U$$1584/A U$$1620/B VGND VGND VPWR VPWR U$$1584/X sky130_fd_sc_hd__xor2_1
XFILLER_203_580 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1595 U$$88/A1 U$$1607/A2 U$$90/A1 U$$1607/B2 VGND VGND VPWR VPWR U$$1596/A sky130_fd_sc_hd__a22o_1
XFILLER_33_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_487 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_79_5 U$$3091/X U$$3224/X U$$3357/X VGND VGND VPWR VPWR dadda_fa_2_80_2/A
+ dadda_fa_2_79_5/A sky130_fd_sc_hd__fa_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$203 final_adder.U$$202/B final_adder.U$$973/B1 final_adder.U$$203/B1
+ VGND VGND VPWR VPWR final_adder.U$$203/X sky130_fd_sc_hd__a21o_1
XTAP_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$214 final_adder.U$$214/A final_adder.U$$214/B VGND VGND VPWR VPWR
+ final_adder.U$$342/B sky130_fd_sc_hd__and2_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$225 final_adder.U$$224/B final_adder.U$$995/B1 final_adder.U$$225/B1
+ VGND VGND VPWR VPWR final_adder.U$$225/X sky130_fd_sc_hd__a21o_1
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$236 final_adder.U$$236/A final_adder.U$$236/B VGND VGND VPWR VPWR
+ final_adder.U$$364/B sky130_fd_sc_hd__and2_1
Xrepeater440 U$$42/A2 VGND VGND VPWR VPWR U$$8/A2 sky130_fd_sc_hd__buf_4
XTAP_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$247 final_adder.U$$9/SUM final_adder.U$$8/COUT final_adder.U$$9/COUT
+ VGND VGND VPWR VPWR final_adder.U$$247/X sky130_fd_sc_hd__a21o_1
XTAP_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater451 U$$4107/A2 VGND VGND VPWR VPWR U$$4103/A2 sky130_fd_sc_hd__buf_4
XFILLER_57_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$258 final_adder.U$$260/B final_adder.U$$258/B VGND VGND VPWR VPWR
+ final_adder.U$$384/B sky130_fd_sc_hd__and2_1
XTAP_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater462 U$$3840/X VGND VGND VPWR VPWR U$$3968/A2 sky130_fd_sc_hd__buf_8
XFILLER_211_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$269 final_adder.U$$268/B final_adder.U$$143/X final_adder.U$$141/X
+ VGND VGND VPWR VPWR final_adder.U$$269/X sky130_fd_sc_hd__a21o_1
XU$$108 U$$654/B1 U$$122/A2 U$$521/A1 U$$122/B2 VGND VGND VPWR VPWR U$$109/A sky130_fd_sc_hd__a22o_1
Xrepeater473 U$$3644/A2 VGND VGND VPWR VPWR U$$3660/A2 sky130_fd_sc_hd__buf_6
Xrepeater484 U$$3517/A2 VGND VGND VPWR VPWR U$$3559/A2 sky130_fd_sc_hd__buf_4
XU$$119 U$$119/A U$$127/B VGND VGND VPWR VPWR U$$119/X sky130_fd_sc_hd__xor2_1
XFILLER_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater495 U$$3255/A2 VGND VGND VPWR VPWR U$$3263/A2 sky130_fd_sc_hd__buf_4
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_482 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4475_1814 VGND VGND VPWR VPWR U$$4475_1814/HI U$$4475/B sky130_fd_sc_hd__conb_1
XFILLER_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_498 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_110_1 U$$3552/X U$$3685/X U$$3818/X VGND VGND VPWR VPWR dadda_fa_4_111_1/A
+ dadda_fa_4_110_2/A sky130_fd_sc_hd__fa_1
Xrepeater1008 U$$2202/B1 VGND VGND VPWR VPWR U$$12/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_111_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1019 U$$3078/B1 VGND VGND VPWR VPWR U$$888/A1 sky130_fd_sc_hd__buf_4
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_863 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_103_0 U$$3937/X U$$4070/X U$$4203/X VGND VGND VPWR VPWR dadda_fa_4_104_0/B
+ dadda_fa_4_103_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_68_5 U$$2271/X U$$2404/X VGND VGND VPWR VPWR dadda_fa_1_69_7/B dadda_fa_2_68_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_972 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput210 c[58] VGND VGND VPWR VPWR input210/X sky130_fd_sc_hd__buf_2
Xinput221 c[68] VGND VGND VPWR VPWR input221/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput232 c[78] VGND VGND VPWR VPWR input232/X sky130_fd_sc_hd__buf_2
Xdadda_fa_3_51_3 dadda_fa_3_51_3/A dadda_fa_3_51_3/B dadda_fa_3_51_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_52_1/B dadda_fa_4_51_2/CIN sky130_fd_sc_hd__fa_1
Xinput243 c[88] VGND VGND VPWR VPWR input243/X sky130_fd_sc_hd__clkbuf_2
XTAP_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_67_3 U$$1338/X U$$1471/X U$$1604/X VGND VGND VPWR VPWR dadda_fa_1_68_6/B
+ dadda_fa_1_67_8/B sky130_fd_sc_hd__fa_1
Xinput254 c[98] VGND VGND VPWR VPWR input254/X sky130_fd_sc_hd__buf_4
XTAP_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_44_2 dadda_fa_3_44_2/A dadda_fa_3_44_2/B dadda_fa_3_44_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_1/A dadda_fa_4_44_2/B sky130_fd_sc_hd__fa_1
XTAP_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$770 final_adder.U$$770/A final_adder.U$$770/B VGND VGND VPWR VPWR
+ final_adder.U$$770/X sky130_fd_sc_hd__and2_1
XTAP_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$781 final_adder.U$$780/B final_adder.U$$701/X final_adder.U$$669/X
+ VGND VGND VPWR VPWR final_adder.U$$781/X sky130_fd_sc_hd__a21o_1
XTAP_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$620 U$$757/A1 U$$624/A2 U$$896/A1 U$$624/B2 VGND VGND VPWR VPWR U$$621/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_37_1 dadda_fa_3_37_1/A dadda_fa_3_37_1/B dadda_fa_3_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_0/CIN dadda_fa_4_37_2/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$792 final_adder.U$$792/A final_adder.U$$792/B VGND VGND VPWR VPWR
+ final_adder.U$$792/X sky130_fd_sc_hd__and2_1
XU$$631 U$$631/A U$$673/B VGND VGND VPWR VPWR U$$631/X sky130_fd_sc_hd__xor2_1
XFILLER_17_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_14_0 dadda_fa_6_14_0/A dadda_fa_6_14_0/B dadda_fa_6_14_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_15_0/B dadda_fa_7_14_0/CIN sky130_fd_sc_hd__fa_1
XU$$642 U$$914/B1 U$$652/A2 U$$918/A1 U$$652/B2 VGND VGND VPWR VPWR U$$643/A sky130_fd_sc_hd__a22o_1
XFILLER_84_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_1032 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$653 U$$653/A U$$684/A VGND VGND VPWR VPWR U$$653/X sky130_fd_sc_hd__xor2_1
XU$$664 U$$938/A1 U$$672/A2 U$$940/A1 U$$668/B2 VGND VGND VPWR VPWR U$$665/A sky130_fd_sc_hd__a22o_1
XU$$675 U$$675/A U$$683/B VGND VGND VPWR VPWR U$$675/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$686 input2/X VGND VGND VPWR VPWR U$$688/B sky130_fd_sc_hd__inv_1
XFILLER_210_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$697 U$$969/B1 U$$711/A2 U$$836/A1 U$$711/B2 VGND VGND VPWR VPWR U$$698/A sky130_fd_sc_hd__a22o_1
XFILLER_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1520 input121/X VGND VGND VPWR VPWR U$$4099/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_96_5 U$$4455/X input252/X dadda_fa_2_96_5/CIN VGND VGND VPWR VPWR dadda_fa_3_97_2/A
+ dadda_fa_4_96_0/A sky130_fd_sc_hd__fa_2
Xrepeater1531 U$$51/B VGND VGND VPWR VPWR U$$43/B sky130_fd_sc_hd__buf_6
Xrepeater1542 U$$4510/A1 VGND VGND VPWR VPWR U$$948/A1 sky130_fd_sc_hd__clkbuf_8
Xrepeater1553 input118/X VGND VGND VPWR VPWR U$$3960/A1 sky130_fd_sc_hd__buf_4
Xrepeater1564 U$$3545/A1 VGND VGND VPWR VPWR U$$118/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_89_4 dadda_fa_2_89_4/A dadda_fa_2_89_4/B dadda_fa_2_89_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_90_1/CIN dadda_fa_3_89_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1575 U$$4502/A1 VGND VGND VPWR VPWR U$$2445/B1 sky130_fd_sc_hd__buf_4
XFILLER_98_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1586 input114/X VGND VGND VPWR VPWR U$$4361/B1 sky130_fd_sc_hd__buf_6
XFILLER_4_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1597 U$$2715/A1 VGND VGND VPWR VPWR U$$932/B1 sky130_fd_sc_hd__buf_6
XFILLER_154_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _327_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_931 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_32_0 U$$71/X U$$204/X U$$337/X VGND VGND VPWR VPWR dadda_fa_3_33_0/B dadda_fa_3_32_2/B
+ sky130_fd_sc_hd__fa_1
XFILLER_78_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2060 U$$2058/B input22/X input24/X U$$2055/Y VGND VGND VPWR VPWR U$$2060/X sky130_fd_sc_hd__a22o_2
XU$$2071 U$$2206/B1 U$$2099/A2 U$$3032/A1 U$$2099/B2 VGND VGND VPWR VPWR U$$2072/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2082 U$$2082/A U$$2092/B VGND VGND VPWR VPWR U$$2082/X sky130_fd_sc_hd__xor2_1
XFILLER_74_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2093 U$$4422/A1 U$$2093/A2 U$$997/B1 U$$2093/B2 VGND VGND VPWR VPWR U$$2094/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1370 U$$1370/A VGND VGND VPWR VPWR U$$1370/Y sky130_fd_sc_hd__inv_1
XFILLER_206_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1381 U$$1381/A U$$1405/B VGND VGND VPWR VPWR U$$1381/X sky130_fd_sc_hd__xor2_1
XFILLER_200_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1392 U$$1666/A1 U$$1422/A2 U$$1666/B1 U$$1422/B2 VGND VGND VPWR VPWR U$$1393/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_119_0 input150/X dadda_fa_5_119_0/B dadda_fa_5_119_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_6_120_0/A dadda_fa_6_119_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1064 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_84_3 U$$2569/X U$$2702/X U$$2835/X VGND VGND VPWR VPWR dadda_fa_2_85_3/A
+ dadda_fa_2_84_5/A sky130_fd_sc_hd__fa_1
XFILLER_171_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_61_2 dadda_fa_4_61_2/A dadda_fa_4_61_2/B dadda_fa_4_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_62_0/CIN dadda_fa_5_61_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_77_2 U$$2156/X U$$2289/X U$$2422/X VGND VGND VPWR VPWR dadda_fa_2_78_1/A
+ dadda_fa_2_77_4/A sky130_fd_sc_hd__fa_1
XFILLER_58_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_54_1 dadda_fa_4_54_1/A dadda_fa_4_54_1/B dadda_fa_4_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/B dadda_fa_5_54_1/B sky130_fd_sc_hd__fa_1
XTAP_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_31_0 dadda_fa_7_31_0/A dadda_fa_7_31_0/B dadda_fa_7_31_0/CIN VGND VGND
+ VPWR VPWR _328_/D _199_/D sky130_fd_sc_hd__fa_2
XFILLER_97_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_47_0 dadda_fa_4_47_0/A dadda_fa_4_47_0/B dadda_fa_4_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/A dadda_fa_5_47_1/A sky130_fd_sc_hd__fa_1
XFILLER_57_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_636 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_371_ _373_/CLK _371_/D VGND VGND VPWR VPWR _371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_99_3 dadda_fa_3_99_3/A dadda_fa_3_99_3/B dadda_fa_3_99_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_100_1/B dadda_fa_4_99_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_72_1 U$$949/X U$$1082/X U$$1215/X VGND VGND VPWR VPWR dadda_fa_1_73_7/B
+ dadda_fa_1_72_8/B sky130_fd_sc_hd__fa_1
XFILLER_89_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_65_0 U$$136/A U$$270/X U$$403/X VGND VGND VPWR VPWR dadda_fa_1_66_5/B
+ dadda_fa_1_65_7/B sky130_fd_sc_hd__fa_1
XFILLER_209_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$450 U$$450/A U$$474/B VGND VGND VPWR VPWR U$$450/X sky130_fd_sc_hd__xor2_1
XFILLER_45_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$461 U$$461/A1 U$$491/A2 U$$461/B1 U$$491/B2 VGND VGND VPWR VPWR U$$462/A sky130_fd_sc_hd__a22o_1
XFILLER_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$472 U$$472/A U$$504/B VGND VGND VPWR VPWR U$$472/X sky130_fd_sc_hd__xor2_1
XU$$483 U$$757/A1 U$$483/A2 U$$483/B1 U$$483/B2 VGND VGND VPWR VPWR U$$484/A sky130_fd_sc_hd__a22o_1
XFILLER_204_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$494 U$$494/A U$$536/B VGND VGND VPWR VPWR U$$494/X sky130_fd_sc_hd__xor2_1
XFILLER_32_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_94_2 U$$3520/X U$$3653/X U$$3786/X VGND VGND VPWR VPWR dadda_fa_3_95_1/A
+ dadda_fa_3_94_3/A sky130_fd_sc_hd__fa_1
XFILLER_99_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1350 U$$184/B VGND VGND VPWR VPWR U$$160/B sky130_fd_sc_hd__buf_4
Xdadda_fa_5_71_1 dadda_fa_5_71_1/A dadda_fa_5_71_1/B dadda_fa_5_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_72_0/B dadda_fa_7_71_0/A sky130_fd_sc_hd__fa_1
Xrepeater1361 U$$2739/A VGND VGND VPWR VPWR U$$2736/B sky130_fd_sc_hd__buf_6
Xdadda_fa_2_87_1 U$$4038/X U$$4171/X U$$4304/X VGND VGND VPWR VPWR dadda_fa_3_88_0/CIN
+ dadda_fa_3_87_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater1372 U$$2569/B VGND VGND VPWR VPWR U$$2577/B sky130_fd_sc_hd__buf_12
XFILLER_119_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1383 input3/X VGND VGND VPWR VPWR U$$808/B sky130_fd_sc_hd__buf_4
XFILLER_113_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_64_0 dadda_fa_5_64_0/A dadda_fa_5_64_0/B dadda_fa_5_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_65_0/A dadda_fa_6_64_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1394 U$$2303/B VGND VGND VPWR VPWR U$$2253/B sky130_fd_sc_hd__buf_6
XFILLER_119_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_63_8 dadda_fa_1_63_8/A dadda_fa_1_63_8/B dadda_fa_1_63_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_64_3/A dadda_fa_3_63_0/A sky130_fd_sc_hd__fa_2
XFILLER_45_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_56_7 U$$3927/B input208/X dadda_fa_1_56_7/CIN VGND VGND VPWR VPWR dadda_fa_2_57_2/CIN
+ dadda_fa_2_56_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_49_6 U$$2499/X U$$2632/X U$$2765/X VGND VGND VPWR VPWR dadda_fa_2_50_2/CIN
+ dadda_fa_2_49_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_199_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_706 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1060 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_90_3 U$$2980/X U$$3113/X VGND VGND VPWR VPWR dadda_fa_2_91_5/A dadda_fa_3_90_0/A
+ sky130_fd_sc_hd__ha_2
XFILLER_210_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_79_0 dadda_fa_7_79_0/A dadda_fa_7_79_0/B dadda_fa_7_79_0/CIN VGND VGND
+ VPWR VPWR _376_/D _247_/D sky130_fd_sc_hd__fa_1
XFILLER_3_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_82_0 dadda_fa_1_82_0/A U$$1368/X U$$1501/X VGND VGND VPWR VPWR dadda_fa_2_83_1/B
+ dadda_fa_2_82_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4209 U$$4209/A U$$4211/B VGND VGND VPWR VPWR U$$4209/X sky130_fd_sc_hd__xor2_1
XFILLER_59_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3508 U$$3508/A U$$3510/B VGND VGND VPWR VPWR U$$3508/X sky130_fd_sc_hd__xor2_1
XFILLER_85_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3519 U$$4478/A1 U$$3549/A2 U$$4478/B1 U$$3549/B2 VGND VGND VPWR VPWR U$$3520/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2807 U$$2807/A U$$2825/B VGND VGND VPWR VPWR U$$2807/X sky130_fd_sc_hd__xor2_1
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2818 U$$4323/B1 U$$2858/A2 U$$4188/B1 U$$2858/B2 VGND VGND VPWR VPWR U$$2819/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_101 _346_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2829 U$$2829/A U$$2845/B VGND VGND VPWR VPWR U$$2829/X sky130_fd_sc_hd__xor2_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 U$$50/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_145 U$$1746/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_156 U$$2149/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_167 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_382 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_423_ _423_/CLK _423_/D VGND VGND VPWR VPWR _423_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_178 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_21 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _198_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_354_ _355_/CLK _354_/D VGND VGND VPWR VPWR _354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_285_ _414_/CLK _285_/D VGND VGND VPWR VPWR _285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_81_0 dadda_fa_6_81_0/A dadda_fa_6_81_0/B dadda_fa_6_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_82_0/B dadda_fa_7_81_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_97_0 dadda_fa_3_97_0/A dadda_fa_3_97_0/B dadda_fa_3_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_0/B dadda_fa_4_97_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_983 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_59_5 dadda_fa_2_59_5/A dadda_fa_2_59_5/B dadda_fa_2_59_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_60_2/A dadda_fa_4_59_0/A sky130_fd_sc_hd__fa_2
XTAP_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 a[15] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_4
XTAP_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$280 U$$280/A1 U$$316/A2 U$$8/A1 U$$316/B2 VGND VGND VPWR VPWR U$$281/A sky130_fd_sc_hd__a22o_1
XFILLER_91_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_472 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$291 U$$291/A U$$379/B VGND VGND VPWR VPWR U$$291/X sky130_fd_sc_hd__xor2_1
XFILLER_162_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$5 _301_/Q _173_/Q VGND VGND VPWR VPWR final_adder.U$$5/COUT final_adder.U$$5/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_173_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput300 output300/A VGND VGND VPWR VPWR o[23] sky130_fd_sc_hd__buf_2
XFILLER_105_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput311 output311/A VGND VGND VPWR VPWR o[33] sky130_fd_sc_hd__buf_2
Xoutput322 output322/A VGND VGND VPWR VPWR o[43] sky130_fd_sc_hd__buf_2
XFILLER_105_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput333 output333/A VGND VGND VPWR VPWR o[53] sky130_fd_sc_hd__buf_2
XFILLER_133_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput344 output344/A VGND VGND VPWR VPWR o[63] sky130_fd_sc_hd__buf_2
Xoutput355 output355/A VGND VGND VPWR VPWR o[73] sky130_fd_sc_hd__buf_2
XFILLER_82_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1180 U$$850/B1 VGND VGND VPWR VPWR U$$987/B1 sky130_fd_sc_hd__buf_4
Xoutput366 output366/A VGND VGND VPWR VPWR o[83] sky130_fd_sc_hd__buf_2
XFILLER_82_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput377 output377/A VGND VGND VPWR VPWR o[93] sky130_fd_sc_hd__buf_2
Xrepeater1191 U$$3453/A1 VGND VGND VPWR VPWR U$$2220/A1 sky130_fd_sc_hd__buf_4
XFILLER_59_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_61_5 U$$3986/X U$$4119/X input214/X VGND VGND VPWR VPWR dadda_fa_2_62_2/A
+ dadda_fa_2_61_5/A sky130_fd_sc_hd__fa_1
XFILLER_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_4 U$$2376/X U$$2509/X U$$2642/X VGND VGND VPWR VPWR dadda_fa_2_55_1/CIN
+ dadda_fa_2_54_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_47_3 U$$1298/X U$$1431/X U$$1564/X VGND VGND VPWR VPWR dadda_fa_2_48_2/B
+ dadda_fa_2_47_5/A sky130_fd_sc_hd__fa_1
XFILLER_82_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_24_2 dadda_fa_4_24_2/A dadda_fa_4_24_2/B dadda_fa_4_24_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_25_0/CIN dadda_fa_5_24_1/CIN sky130_fd_sc_hd__fa_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_17_1 U$$1105/X input165/X dadda_fa_4_17_1/CIN VGND VGND VPWR VPWR dadda_fa_5_18_0/B
+ dadda_fa_5_17_1/B sky130_fd_sc_hd__fa_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4006 U$$4006/A U$$4044/B VGND VGND VPWR VPWR U$$4006/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_20_3 U$$1244/X U$$1377/X VGND VGND VPWR VPWR dadda_fa_4_21_1/B dadda_ha_3_20_3/SUM
+ sky130_fd_sc_hd__ha_1
XU$$4017 input74/X U$$4107/A2 U$$4019/A1 U$$4107/B2 VGND VGND VPWR VPWR U$$4018/A
+ sky130_fd_sc_hd__a22o_1
XU$$4028 U$$4028/A U$$4044/B VGND VGND VPWR VPWR U$$4028/X sky130_fd_sc_hd__xor2_1
XFILLER_115_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4039 U$$4176/A1 U$$3977/X U$$4176/B1 U$$3978/X VGND VGND VPWR VPWR U$$4040/A sky130_fd_sc_hd__a22o_1
XFILLER_111_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3305 U$$3305/A U$$3395/B VGND VGND VPWR VPWR U$$3305/X sky130_fd_sc_hd__xor2_1
XFILLER_150_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3316 U$$4410/B1 U$$3320/A2 U$$989/A1 U$$3320/B2 VGND VGND VPWR VPWR U$$3317/A
+ sky130_fd_sc_hd__a22o_1
XU$$3327 U$$3327/A U$$3349/B VGND VGND VPWR VPWR U$$3327/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3338 U$$4434/A1 U$$3292/X U$$4297/B1 U$$3293/X VGND VGND VPWR VPWR U$$3339/A sky130_fd_sc_hd__a22o_1
XU$$2604 input32/X VGND VGND VPWR VPWR U$$2606/B sky130_fd_sc_hd__inv_1
XU$$3349 U$$3349/A U$$3349/B VGND VGND VPWR VPWR U$$3349/X sky130_fd_sc_hd__xor2_1
XU$$2615 U$$3026/A1 U$$2625/A2 U$$3028/A1 U$$2625/B2 VGND VGND VPWR VPWR U$$2616/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2626 U$$2626/A U$$2658/B VGND VGND VPWR VPWR U$$2626/X sky130_fd_sc_hd__xor2_1
XFILLER_46_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2637 U$$32/B1 U$$2727/A2 U$$4146/A1 U$$2727/B2 VGND VGND VPWR VPWR U$$2638/A sky130_fd_sc_hd__a22o_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2648 U$$2648/A U$$2736/B VGND VGND VPWR VPWR U$$2648/X sky130_fd_sc_hd__xor2_1
XU$$1903 U$$2312/B1 U$$1785/X U$$2316/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1904/A
+ sky130_fd_sc_hd__a22o_1
XU$$2659 U$$3344/A1 U$$2691/A2 U$$58/A1 U$$2691/B2 VGND VGND VPWR VPWR U$$2660/A sky130_fd_sc_hd__a22o_1
XFILLER_61_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1914 U$$1914/A U$$1914/B VGND VGND VPWR VPWR U$$1914/X sky130_fd_sc_hd__xor2_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1925 U$$1925/A U$$1993/B VGND VGND VPWR VPWR U$$1925/X sky130_fd_sc_hd__xor2_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1936 U$$3032/A1 U$$1970/A2 U$$979/A1 U$$1970/B2 VGND VGND VPWR VPWR U$$1937/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1947 U$$1947/A U$$2009/B VGND VGND VPWR VPWR U$$1947/X sky130_fd_sc_hd__xor2_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1958 U$$860/B1 U$$2022/A2 U$$727/A1 U$$2022/B2 VGND VGND VPWR VPWR U$$1959/A sky130_fd_sc_hd__a22o_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_406_ _407_/CLK _406_/D VGND VGND VPWR VPWR _406_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1969 U$$1969/A U$$1971/B VGND VGND VPWR VPWR U$$1969/X sky130_fd_sc_hd__xor2_1
XFILLER_203_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_337_ _337_/CLK _337_/D VGND VGND VPWR VPWR _337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_338 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_268_ _397_/CLK _268_/D VGND VGND VPWR VPWR _268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_199_ _327_/CLK _199_/D VGND VGND VPWR VPWR _199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_71_4 dadda_fa_2_71_4/A dadda_fa_2_71_4/B dadda_fa_2_71_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_1/CIN dadda_fa_3_71_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_64_3 dadda_fa_2_64_3/A dadda_fa_2_64_3/B dadda_fa_2_64_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/B dadda_fa_3_64_3/B sky130_fd_sc_hd__fa_1
Xrepeater803 U$$2459/B2 VGND VGND VPWR VPWR U$$2463/B2 sky130_fd_sc_hd__buf_4
XFILLER_57_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater814 U$$2091/B2 VGND VGND VPWR VPWR U$$2093/B2 sky130_fd_sc_hd__buf_4
XFILLER_38_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater825 U$$2022/B2 VGND VGND VPWR VPWR U$$2016/B2 sky130_fd_sc_hd__buf_6
XFILLER_96_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_57_2 dadda_fa_2_57_2/A dadda_fa_2_57_2/B dadda_fa_2_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/A dadda_fa_3_57_3/A sky130_fd_sc_hd__fa_1
Xrepeater836 U$$1786/X VGND VGND VPWR VPWR U$$1903/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_110_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater847 U$$1621/B2 VGND VGND VPWR VPWR U$$1575/B2 sky130_fd_sc_hd__buf_4
Xrepeater858 U$$259/B2 VGND VGND VPWR VPWR U$$209/B2 sky130_fd_sc_hd__buf_4
XU$$10 U$$8/B1 U$$8/A2 U$$12/A1 U$$8/B2 VGND VGND VPWR VPWR U$$11/A sky130_fd_sc_hd__a22o_1
Xrepeater869 U$$1375/X VGND VGND VPWR VPWR U$$1470/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_34_1 dadda_fa_5_34_1/A dadda_fa_5_34_1/B dadda_fa_5_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_35_0/B dadda_fa_7_34_0/A sky130_fd_sc_hd__fa_1
XU$$21 U$$21/A U$$43/B VGND VGND VPWR VPWR U$$21/X sky130_fd_sc_hd__xor2_1
XU$$32 U$$32/A1 U$$50/A2 U$$32/B1 U$$50/B2 VGND VGND VPWR VPWR U$$33/A sky130_fd_sc_hd__a22o_1
XU$$43 U$$43/A U$$43/B VGND VGND VPWR VPWR U$$43/X sky130_fd_sc_hd__xor2_1
XFILLER_37_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_27_0 dadda_fa_5_27_0/A dadda_fa_5_27_0/B dadda_fa_5_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_28_0/A dadda_fa_6_27_0/CIN sky130_fd_sc_hd__fa_1
XU$$54 U$$54/A1 U$$98/A2 U$$56/A1 U$$98/B2 VGND VGND VPWR VPWR U$$55/A sky130_fd_sc_hd__a22o_1
XU$$3850 input98/X U$$3878/A2 U$$3852/A1 U$$3878/B2 VGND VGND VPWR VPWR U$$3851/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$65 U$$65/A U$$85/B VGND VGND VPWR VPWR U$$65/X sky130_fd_sc_hd__xor2_1
XU$$3861 U$$3861/A U$$3875/B VGND VGND VPWR VPWR U$$3861/X sky130_fd_sc_hd__xor2_1
XFILLER_65_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$76 U$$76/A1 U$$80/A2 U$$78/A1 U$$80/B2 VGND VGND VPWR VPWR U$$77/A sky130_fd_sc_hd__a22o_1
XU$$87 U$$87/A U$$99/B VGND VGND VPWR VPWR U$$87/X sky130_fd_sc_hd__xor2_1
XU$$3872 U$$4009/A1 U$$3874/A2 U$$4422/A1 U$$3874/B2 VGND VGND VPWR VPWR U$$3873/A
+ sky130_fd_sc_hd__a22o_1
XU$$3883 U$$3883/A U$$3927/B VGND VGND VPWR VPWR U$$3883/X sky130_fd_sc_hd__xor2_1
XU$$98 U$$98/A1 U$$98/A2 U$$98/B1 U$$98/B2 VGND VGND VPWR VPWR U$$99/A sky130_fd_sc_hd__a22o_1
XU$$3894 U$$4442/A1 U$$3840/X input83/X U$$3841/X VGND VGND VPWR VPWR U$$3895/A sky130_fd_sc_hd__a22o_1
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_12 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_23 _337_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_34 _339_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_56 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 _342_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_78 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 _344_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_101_0 dadda_fa_5_101_0/A dadda_fa_5_101_0/B dadda_fa_5_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_102_0/A dadda_fa_6_101_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_146_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_52_1 U$$776/X U$$909/X U$$1042/X VGND VGND VPWR VPWR dadda_fa_2_53_0/CIN
+ dadda_fa_2_52_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_45_0 U$$97/X U$$230/X U$$363/X VGND VGND VPWR VPWR dadda_fa_2_46_2/A dadda_fa_2_45_4/B
+ sky130_fd_sc_hd__fa_1
XFILLER_83_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_920 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_986 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_327 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1015 final_adder.U$$244/A final_adder.U$$625/X final_adder.U$$245/A2
+ VGND VGND VPWR VPWR final_adder.U$$1035/B sky130_fd_sc_hd__a21o_1
XFILLER_7_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1026 final_adder.U$$252/A final_adder.U$$255/X VGND VGND VPWR VPWR
+ output307/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1037 final_adder.U$$242/B final_adder.U$$1037/B VGND VGND VPWR VPWR
+ output289/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1048 final_adder.U$$230/A final_adder.U$$731/X VGND VGND VPWR VPWR
+ output301/A sky130_fd_sc_hd__xor2_1
XFILLER_194_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$1059 final_adder.U$$220/B final_adder.U$$991/X VGND VGND VPWR VPWR
+ output313/A sky130_fd_sc_hd__xor2_1
XFILLER_164_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_81_3 dadda_fa_3_81_3/A dadda_fa_3_81_3/B dadda_fa_3_81_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_82_1/B dadda_fa_4_81_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_180_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_74_2 dadda_fa_3_74_2/A dadda_fa_3_74_2/B dadda_fa_3_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_1/A dadda_fa_4_74_2/B sky130_fd_sc_hd__fa_1
XFILLER_127_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_67_1 dadda_fa_3_67_1/A dadda_fa_3_67_1/B dadda_fa_3_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_0/CIN dadda_fa_4_67_2/A sky130_fd_sc_hd__fa_1
XFILLER_26_1238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_44_0 dadda_fa_6_44_0/A dadda_fa_6_44_0/B dadda_fa_6_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_45_0/B dadda_fa_7_44_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3102 U$$3376/A1 U$$3108/A2 U$$3102/B1 U$$3108/B2 VGND VGND VPWR VPWR U$$3103/A
+ sky130_fd_sc_hd__a22o_1
XU$$3113 U$$3113/A U$$3151/A VGND VGND VPWR VPWR U$$3113/X sky130_fd_sc_hd__xor2_1
XFILLER_93_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3124 U$$384/A1 U$$3124/A2 U$$3946/B1 U$$3124/B2 VGND VGND VPWR VPWR U$$3125/A
+ sky130_fd_sc_hd__a22o_1
XU$$3135 U$$3135/A U$$3150/A VGND VGND VPWR VPWR U$$3135/X sky130_fd_sc_hd__xor2_1
XU$$3146 U$$3281/B1 U$$3148/A2 U$$3148/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3147/A
+ sky130_fd_sc_hd__a22o_1
XU$$2401 U$$4043/B1 U$$2333/X U$$3499/A1 U$$2334/X VGND VGND VPWR VPWR U$$2402/A sky130_fd_sc_hd__a22o_1
XU$$3157 U$$3157/A1 U$$3207/A2 U$$3159/A1 U$$3207/B2 VGND VGND VPWR VPWR U$$3158/A
+ sky130_fd_sc_hd__a22o_1
XU$$2412 U$$2412/A U$$2446/B VGND VGND VPWR VPWR U$$2412/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_103_2 dadda_fa_4_103_2/A dadda_fa_4_103_2/B dadda_fa_4_103_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_104_0/CIN dadda_fa_5_103_1/CIN sky130_fd_sc_hd__fa_1
XU$$3168 U$$3168/A U$$3188/B VGND VGND VPWR VPWR U$$3168/X sky130_fd_sc_hd__xor2_1
XU$$2423 U$$3245/A1 U$$2449/A2 U$$3245/B1 U$$2449/B2 VGND VGND VPWR VPWR U$$2424/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2434 U$$2434/A U$$2446/B VGND VGND VPWR VPWR U$$2434/X sky130_fd_sc_hd__xor2_1
XU$$3179 input66/X U$$3229/A2 input67/X U$$3227/B2 VGND VGND VPWR VPWR U$$3180/A sky130_fd_sc_hd__a22o_1
XU$$2445 U$$936/B1 U$$2449/A2 U$$2445/B1 U$$2449/B2 VGND VGND VPWR VPWR U$$2446/A
+ sky130_fd_sc_hd__a22o_1
XU$$1700 U$$741/A1 U$$1706/A2 U$$878/B1 U$$1706/B2 VGND VGND VPWR VPWR U$$1701/A sky130_fd_sc_hd__a22o_1
XFILLER_146_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1711 U$$1711/A U$$1721/B VGND VGND VPWR VPWR U$$1711/X sky130_fd_sc_hd__xor2_1
XU$$2456 U$$2456/A U$$2465/A VGND VGND VPWR VPWR U$$2456/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_94_0_1859 VGND VGND VPWR VPWR dadda_fa_1_94_0/A dadda_fa_1_94_0_1859/LO
+ sky130_fd_sc_hd__conb_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2467 input30/X VGND VGND VPWR VPWR U$$2469/B sky130_fd_sc_hd__inv_1
XU$$1722 U$$78/A1 U$$1750/A2 U$$80/A1 U$$1750/B2 VGND VGND VPWR VPWR U$$1723/A sky130_fd_sc_hd__a22o_1
XFILLER_188_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1733 U$$1733/A U$$1779/B VGND VGND VPWR VPWR U$$1733/X sky130_fd_sc_hd__xor2_1
XU$$2478 U$$3026/A1 U$$2524/A2 U$$3028/A1 U$$2524/B2 VGND VGND VPWR VPWR U$$2479/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2489 U$$2489/A U$$2491/B VGND VGND VPWR VPWR U$$2489/X sky130_fd_sc_hd__xor2_1
XU$$1744 U$$2701/B1 U$$1770/A2 U$$2292/B1 U$$1770/B2 VGND VGND VPWR VPWR U$$1745/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1755 U$$1755/A U$$1765/B VGND VGND VPWR VPWR U$$1755/X sky130_fd_sc_hd__xor2_1
XFILLER_61_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1766 U$$2312/B1 U$$1770/A2 U$$2316/A1 U$$1770/B2 VGND VGND VPWR VPWR U$$1767/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1777 U$$1777/A U$$1779/B VGND VGND VPWR VPWR U$$1777/X sky130_fd_sc_hd__xor2_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1788 U$$1788/A U$$1820/B VGND VGND VPWR VPWR U$$1788/X sky130_fd_sc_hd__xor2_1
XFILLER_72_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1799 U$$1799/A1 U$$1831/A2 U$$1799/B1 U$$1831/B2 VGND VGND VPWR VPWR U$$1800/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_117_0 dadda_fa_7_117_0/A dadda_fa_7_117_0/B dadda_fa_7_117_0/CIN VGND
+ VGND VPWR VPWR _414_/D _285_/D sky130_fd_sc_hd__fa_1
XFILLER_30_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 a[18] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_2
Xinput21 a[28] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_1
Xinput32 a[38] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput43 a[48] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
Xinput54 a[58] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_1
Xinput65 b[0] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__buf_8
XFILLER_116_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput76 b[1] VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__buf_8
Xinput87 b[2] VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__buf_6
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput98 b[3] VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__buf_8
XFILLER_192_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater600 U$$1621/A2 VGND VGND VPWR VPWR U$$1575/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_62_0 dadda_fa_2_62_0/A dadda_fa_2_62_0/B dadda_fa_2_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_0/B dadda_fa_3_62_2/B sky130_fd_sc_hd__fa_1
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$407 final_adder.U$$406/B final_adder.U$$285/X final_adder.U$$281/X
+ VGND VGND VPWR VPWR final_adder.U$$407/X sky130_fd_sc_hd__a21o_1
Xrepeater611 U$$259/A2 VGND VGND VPWR VPWR U$$209/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$418 final_adder.U$$422/B final_adder.U$$418/B VGND VGND VPWR VPWR
+ final_adder.U$$542/B sky130_fd_sc_hd__and2_1
Xrepeater622 U$$1374/X VGND VGND VPWR VPWR U$$1470/A2 sky130_fd_sc_hd__buf_4
XFILLER_97_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$429 final_adder.U$$428/B final_adder.U$$307/X final_adder.U$$303/X
+ VGND VGND VPWR VPWR final_adder.U$$429/X sky130_fd_sc_hd__a21o_1
Xrepeater633 U$$1174/A2 VGND VGND VPWR VPWR U$$1138/A2 sky130_fd_sc_hd__buf_4
Xrepeater644 U$$1057/B2 VGND VGND VPWR VPWR U$$965/B2 sky130_fd_sc_hd__buf_6
XFILLER_85_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater655 U$$783/B2 VGND VGND VPWR VPWR U$$711/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_38_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater666 U$$678/B2 VGND VGND VPWR VPWR U$$652/B2 sky130_fd_sc_hd__buf_4
Xrepeater677 U$$4252/X VGND VGND VPWR VPWR U$$4373/B2 sky130_fd_sc_hd__buf_6
XFILLER_26_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater688 U$$4115/X VGND VGND VPWR VPWR U$$4176/B2 sky130_fd_sc_hd__buf_4
XFILLER_203_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater699 U$$4107/B2 VGND VGND VPWR VPWR U$$4043/B2 sky130_fd_sc_hd__buf_12
XU$$4370 U$$4370/A U$$4370/B VGND VGND VPWR VPWR U$$4370/X sky130_fd_sc_hd__xor2_1
XU$$4381 U$$4516/B1 U$$4381/A2 U$$4381/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4382/A
+ sky130_fd_sc_hd__a22o_1
XU$$4392 U$$4392/A1 U$$4388/X U$$4394/A1 U$$4432/B2 VGND VGND VPWR VPWR U$$4393/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3680 U$$3680/A1 U$$3680/A2 U$$118/B1 U$$3680/B2 VGND VGND VPWR VPWR U$$3681/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3691 U$$3691/A U$$3698/A VGND VGND VPWR VPWR U$$3691/X sky130_fd_sc_hd__xor2_1
XFILLER_53_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_931 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2990 U$$2990/A U$$3013/A VGND VGND VPWR VPWR U$$2990/X sky130_fd_sc_hd__xor2_1
XFILLER_34_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_91_2 dadda_fa_4_91_2/A dadda_fa_4_91_2/B dadda_fa_4_91_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_92_0/CIN dadda_fa_5_91_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_84_1 dadda_fa_4_84_1/A dadda_fa_4_84_1/B dadda_fa_4_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/B dadda_fa_5_84_1/B sky130_fd_sc_hd__fa_1
XFILLER_88_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_61_0 dadda_fa_7_61_0/A dadda_fa_7_61_0/B dadda_fa_7_61_0/CIN VGND VGND
+ VPWR VPWR _358_/D _229_/D sky130_fd_sc_hd__fa_1
XFILLER_164_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_77_0 dadda_fa_4_77_0/A dadda_fa_4_77_0/B dadda_fa_4_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/A dadda_fa_5_77_1/A sky130_fd_sc_hd__fa_1
XFILLER_0_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$941 final_adder.U$$170/A final_adder.U$$879/X final_adder.U$$941/B1
+ VGND VGND VPWR VPWR final_adder.U$$941/X sky130_fd_sc_hd__a21o_1
XFILLER_189_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$963 final_adder.U$$192/A final_adder.U$$805/X final_adder.U$$963/B1
+ VGND VGND VPWR VPWR final_adder.U$$963/X sky130_fd_sc_hd__a21o_1
XFILLER_169_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$802 U$$802/A U$$808/B VGND VGND VPWR VPWR U$$802/X sky130_fd_sc_hd__xor2_1
XFILLER_60_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$813 U$$950/A1 U$$689/X U$$950/B1 U$$690/X VGND VGND VPWR VPWR U$$814/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$985 final_adder.U$$214/A final_adder.U$$827/X final_adder.U$$985/B1
+ VGND VGND VPWR VPWR final_adder.U$$985/X sky130_fd_sc_hd__a21o_1
XU$$824 U$$959/A VGND VGND VPWR VPWR U$$824/Y sky130_fd_sc_hd__inv_1
XU$$835 U$$835/A U$$847/B VGND VGND VPWR VPWR U$$835/X sky130_fd_sc_hd__xor2_1
XFILLER_29_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_73 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$846 U$$983/A1 U$$872/A2 U$$846/B1 U$$872/B2 VGND VGND VPWR VPWR U$$847/A sky130_fd_sc_hd__a22o_1
XU$$857 U$$857/A U$$929/B VGND VGND VPWR VPWR U$$857/X sky130_fd_sc_hd__xor2_1
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1007 U$$3747/A1 U$$1057/A2 U$$2925/B1 U$$1057/B2 VGND VGND VPWR VPWR U$$1008/A
+ sky130_fd_sc_hd__a22o_1
XU$$868 U$$46/A1 U$$872/A2 U$$48/A1 U$$872/B2 VGND VGND VPWR VPWR U$$869/A sky130_fd_sc_hd__a22o_1
XU$$1018 U$$1018/A U$$994/B VGND VGND VPWR VPWR U$$1018/X sky130_fd_sc_hd__xor2_1
XU$$879 U$$879/A U$$883/B VGND VGND VPWR VPWR U$$879/X sky130_fd_sc_hd__xor2_1
XFILLER_204_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1029 U$$892/A1 U$$1083/A2 U$$894/A1 U$$1083/B2 VGND VGND VPWR VPWR U$$1030/A sky130_fd_sc_hd__a22o_1
XFILLER_204_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_794 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1702 input100/X VGND VGND VPWR VPWR U$$912/A1 sky130_fd_sc_hd__buf_4
XFILLER_208_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1076 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_859 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_41_5 dadda_fa_2_41_5/A dadda_fa_2_41_5/B dadda_fa_2_41_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_42_2/A dadda_fa_4_41_0/A sky130_fd_sc_hd__fa_2
XFILLER_47_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2220 U$$2220/A1 U$$2272/A2 U$$2357/B1 U$$2272/B2 VGND VGND VPWR VPWR U$$2221/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_34_4 U$$1937/X U$$2070/X U$$2203/X VGND VGND VPWR VPWR dadda_fa_3_35_1/CIN
+ dadda_fa_3_34_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2231 U$$2231/A U$$2253/B VGND VGND VPWR VPWR U$$2231/X sky130_fd_sc_hd__xor2_1
XU$$2242 U$$3749/A1 U$$2284/A2 U$$3749/B1 U$$2284/B2 VGND VGND VPWR VPWR U$$2243/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2253 U$$2253/A U$$2253/B VGND VGND VPWR VPWR U$$2253/X sky130_fd_sc_hd__xor2_1
XU$$2264 U$$894/A1 U$$2308/A2 U$$3499/A1 U$$2308/B2 VGND VGND VPWR VPWR U$$2265/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1530 U$$1530/A U$$1546/B VGND VGND VPWR VPWR U$$1530/X sky130_fd_sc_hd__xor2_1
XU$$2275 U$$2275/A U$$2303/B VGND VGND VPWR VPWR U$$2275/X sky130_fd_sc_hd__xor2_1
XFILLER_179_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2286 U$$914/B1 U$$2326/A2 U$$918/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2287/A sky130_fd_sc_hd__a22o_1
XFILLER_16_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1541 U$$2363/A1 U$$1591/A2 U$$995/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1542/A
+ sky130_fd_sc_hd__a22o_1
XU$$1552 U$$1552/A U$$1558/B VGND VGND VPWR VPWR U$$1552/X sky130_fd_sc_hd__xor2_1
XU$$2297 U$$2297/A U$$2317/B VGND VGND VPWR VPWR U$$2297/X sky130_fd_sc_hd__xor2_1
XU$$1563 U$$330/A1 U$$1591/A2 U$$56/B1 U$$1591/B2 VGND VGND VPWR VPWR U$$1564/A sky130_fd_sc_hd__a22o_1
XU$$1574 U$$1574/A U$$1574/B VGND VGND VPWR VPWR U$$1574/X sky130_fd_sc_hd__xor2_1
XU$$1585 U$$4323/B1 U$$1621/A2 U$$80/A1 U$$1621/B2 VGND VGND VPWR VPWR U$$1586/A sky130_fd_sc_hd__a22o_1
XFILLER_176_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1596 U$$1596/A U$$1608/B VGND VGND VPWR VPWR U$$1596/X sky130_fd_sc_hd__xor2_1
XFILLER_147_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1066 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1099 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_94_0 dadda_fa_5_94_0/A dadda_fa_5_94_0/B dadda_fa_5_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_95_0/A dadda_fa_6_94_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_79_6 U$$3490/X U$$3623/X U$$3756/X VGND VGND VPWR VPWR dadda_fa_2_80_2/B
+ dadda_fa_2_79_5/B sky130_fd_sc_hd__fa_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$204 final_adder.U$$204/A final_adder.U$$204/B VGND VGND VPWR VPWR
+ final_adder.U$$332/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$215 final_adder.U$$214/B final_adder.U$$985/B1 final_adder.U$$215/B1
+ VGND VGND VPWR VPWR final_adder.U$$215/X sky130_fd_sc_hd__a21o_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_945 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$226 final_adder.U$$226/A final_adder.U$$226/B VGND VGND VPWR VPWR
+ final_adder.U$$354/B sky130_fd_sc_hd__and2_1
XFILLER_170_1187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater430 U$$415/X VGND VGND VPWR VPWR U$$537/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$237 final_adder.U$$236/B final_adder.U$$237/A2 final_adder.U$$237/B1
+ VGND VGND VPWR VPWR final_adder.U$$237/X sky130_fd_sc_hd__a21o_1
Xrepeater441 U$$50/A2 VGND VGND VPWR VPWR U$$42/A2 sky130_fd_sc_hd__buf_2
XTAP_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$248 final_adder.U$$6/SUM final_adder.U$$7/SUM VGND VGND VPWR VPWR
+ final_adder.U$$376/B sky130_fd_sc_hd__and2_1
XTAP_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater452 U$$4107/A2 VGND VGND VPWR VPWR U$$4043/A2 sky130_fd_sc_hd__buf_12
Xfinal_adder.U$$259 final_adder.U$$258/B final_adder.U$$133/X final_adder.U$$131/X
+ VGND VGND VPWR VPWR final_adder.U$$259/X sky130_fd_sc_hd__a21o_1
Xrepeater463 U$$3753/A2 VGND VGND VPWR VPWR U$$3793/A2 sky130_fd_sc_hd__buf_6
XU$$109 U$$109/A U$$111/B VGND VGND VPWR VPWR U$$109/X sky130_fd_sc_hd__xor2_1
Xrepeater474 U$$3686/A2 VGND VGND VPWR VPWR U$$3680/A2 sky130_fd_sc_hd__buf_4
XFILLER_26_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater485 U$$3517/A2 VGND VGND VPWR VPWR U$$3489/A2 sky130_fd_sc_hd__buf_6
Xrepeater496 U$$3285/A2 VGND VGND VPWR VPWR U$$3277/A2 sky130_fd_sc_hd__buf_4
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_951 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1009 U$$2202/B1 VGND VGND VPWR VPWR U$$969/B1 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_110_2 U$$3951/X U$$4084/X U$$4217/X VGND VGND VPWR VPWR dadda_fa_4_111_1/B
+ dadda_fa_4_110_2/B sky130_fd_sc_hd__fa_1
XFILLER_175_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_103_1 U$$4336/X U$$4469/X input133/X VGND VGND VPWR VPWR dadda_fa_4_104_0/CIN
+ dadda_fa_4_103_2/A sky130_fd_sc_hd__fa_1
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_599 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_396 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput200 c[49] VGND VGND VPWR VPWR input200/X sky130_fd_sc_hd__buf_2
Xinput211 c[59] VGND VGND VPWR VPWR input211/X sky130_fd_sc_hd__buf_2
XFILLER_89_984 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput222 c[69] VGND VGND VPWR VPWR input222/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_124_0 dadda_fa_6_124_0/A dadda_fa_6_124_0/B dadda_fa_6_124_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_125_0/B dadda_fa_7_124_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_191_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput233 c[79] VGND VGND VPWR VPWR input233/X sky130_fd_sc_hd__buf_2
XTAP_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput244 c[89] VGND VGND VPWR VPWR input244/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_67_4 U$$1737/X U$$1870/X U$$2003/X VGND VGND VPWR VPWR dadda_fa_1_68_6/CIN
+ dadda_fa_1_67_8/CIN sky130_fd_sc_hd__fa_1
Xinput255 c[99] VGND VGND VPWR VPWR input255/X sky130_fd_sc_hd__buf_4
XFILLER_76_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_44_3 dadda_fa_3_44_3/A dadda_fa_3_44_3/B dadda_fa_3_44_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_45_1/B dadda_fa_4_44_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_208_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$760 final_adder.U$$792/B final_adder.U$$760/B VGND VGND VPWR VPWR
+ final_adder.U$$760/X sky130_fd_sc_hd__and2_1
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$771 final_adder.U$$770/B final_adder.U$$691/X final_adder.U$$659/X
+ VGND VGND VPWR VPWR final_adder.U$$771/X sky130_fd_sc_hd__a21o_1
XTAP_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$610 U$$610/A1 U$$636/A2 U$$610/B1 U$$636/B2 VGND VGND VPWR VPWR U$$611/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$782 final_adder.U$$782/A final_adder.U$$782/B VGND VGND VPWR VPWR
+ final_adder.U$$782/X sky130_fd_sc_hd__and2_1
XTAP_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$621 U$$621/A U$$625/B VGND VGND VPWR VPWR U$$621/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_37_2 dadda_fa_3_37_2/A dadda_fa_3_37_2/B dadda_fa_3_37_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_1/A dadda_fa_4_37_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$793 final_adder.U$$792/B final_adder.U$$713/X final_adder.U$$681/X
+ VGND VGND VPWR VPWR final_adder.U$$793/X sky130_fd_sc_hd__a21o_1
XU$$632 U$$84/A1 U$$636/A2 U$$84/B1 U$$636/B2 VGND VGND VPWR VPWR U$$633/A sky130_fd_sc_hd__a22o_1
XU$$643 U$$643/A U$$651/B VGND VGND VPWR VPWR U$$643/X sky130_fd_sc_hd__xor2_1
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$654 U$$654/A1 U$$678/A2 U$$654/B1 U$$678/B2 VGND VGND VPWR VPWR U$$655/A sky130_fd_sc_hd__a22o_1
XFILLER_1_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$665 U$$665/A U$$673/B VGND VGND VPWR VPWR U$$665/X sky130_fd_sc_hd__xor2_1
XFILLER_182_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$676 U$$676/A1 U$$678/A2 U$$676/B1 U$$678/B2 VGND VGND VPWR VPWR U$$677/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$687 U$$808/B VGND VGND VPWR VPWR U$$687/Y sky130_fd_sc_hd__inv_1
XU$$698 U$$698/A U$$784/B VGND VGND VPWR VPWR U$$698/X sky130_fd_sc_hd__xor2_1
XFILLER_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_551 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1510 U$$3829/A1 VGND VGND VPWR VPWR U$$4375/B1 sky130_fd_sc_hd__buf_4
XFILLER_172_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1521 U$$3032/A1 VGND VGND VPWR VPWR U$$1799/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1532 U$$81/B VGND VGND VPWR VPWR U$$51/B sky130_fd_sc_hd__buf_6
XFILLER_125_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1543 U$$3960/B1 VGND VGND VPWR VPWR U$$4510/A1 sky130_fd_sc_hd__buf_6
Xrepeater1554 input118/X VGND VGND VPWR VPWR U$$3684/B1 sky130_fd_sc_hd__buf_4
Xrepeater1565 input116/X VGND VGND VPWR VPWR U$$3545/A1 sky130_fd_sc_hd__buf_4
XFILLER_4_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_89_5 dadda_fa_2_89_5/A dadda_fa_2_89_5/B dadda_fa_2_89_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_90_2/A dadda_fa_4_89_0/A sky130_fd_sc_hd__fa_2
Xrepeater1576 input115/X VGND VGND VPWR VPWR U$$4502/A1 sky130_fd_sc_hd__buf_4
Xrepeater1587 U$$4498/A1 VGND VGND VPWR VPWR U$$660/B1 sky130_fd_sc_hd__buf_6
Xrepeater1598 U$$2715/A1 VGND VGND VPWR VPWR U$$934/A1 sky130_fd_sc_hd__buf_4
XFILLER_113_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_26_2 U$$857/X U$$990/X VGND VGND VPWR VPWR dadda_fa_3_27_3/A dadda_fa_4_26_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_95_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_32_1 U$$470/X U$$603/X U$$736/X VGND VGND VPWR VPWR dadda_fa_3_33_0/CIN
+ dadda_fa_3_32_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_35_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_25_0 U$$57/X U$$190/X U$$323/X VGND VGND VPWR VPWR dadda_fa_3_26_2/CIN
+ dadda_fa_3_25_3/CIN sky130_fd_sc_hd__fa_1
XU$$2050 U$$4103/B1 U$$2052/A2 U$$4242/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2051/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2061 U$$2061/A1 U$$2093/A2 U$$2198/B1 U$$2093/B2 VGND VGND VPWR VPWR U$$2062/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2072 U$$2072/A U$$2100/B VGND VGND VPWR VPWR U$$2072/X sky130_fd_sc_hd__xor2_1
XU$$2083 U$$2220/A1 U$$2091/A2 U$$2357/B1 U$$2091/B2 VGND VGND VPWR VPWR U$$2084/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_161_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2094 U$$2094/A U$$2094/B VGND VGND VPWR VPWR U$$2094/X sky130_fd_sc_hd__xor2_1
XFILLER_50_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1360 U$$1360/A U$$1366/B VGND VGND VPWR VPWR U$$1360/X sky130_fd_sc_hd__xor2_1
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1371 input13/X VGND VGND VPWR VPWR U$$1373/B sky130_fd_sc_hd__inv_1
XU$$1382 U$$2202/B1 U$$1404/A2 U$$2069/A1 U$$1404/B2 VGND VGND VPWR VPWR U$$1383/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1393 U$$1393/A U$$1423/B VGND VGND VPWR VPWR U$$1393/X sky130_fd_sc_hd__xor2_1
XFILLER_200_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_119_1 dadda_fa_5_119_1/A dadda_fa_5_119_1/B dadda_fa_5_119_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_120_0/B dadda_fa_7_119_0/A sky130_fd_sc_hd__fa_1
XFILLER_164_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1076 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_84_4 U$$2968/X U$$3101/X U$$3234/X VGND VGND VPWR VPWR dadda_fa_2_85_3/B
+ dadda_fa_2_84_5/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_77_3 U$$2555/X U$$2688/X U$$2821/X VGND VGND VPWR VPWR dadda_fa_2_78_1/B
+ dadda_fa_2_77_4/B sky130_fd_sc_hd__fa_1
XFILLER_98_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_54_2 dadda_fa_4_54_2/A dadda_fa_4_54_2/B dadda_fa_4_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_55_0/CIN dadda_fa_5_54_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_47_1 dadda_fa_4_47_1/A dadda_fa_4_47_1/B dadda_fa_4_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/B dadda_fa_5_47_1/B sky130_fd_sc_hd__fa_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_24_0 dadda_fa_7_24_0/A dadda_fa_7_24_0/B dadda_fa_7_24_0/CIN VGND VGND
+ VPWR VPWR _321_/D _192_/D sky130_fd_sc_hd__fa_2
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ _370_/CLK _370_/D VGND VGND VPWR VPWR _370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1048 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1093_1710 VGND VGND VPWR VPWR U$$1093_1710/HI U$$1093/B1 sky130_fd_sc_hd__conb_1
XFILLER_181_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_72_2 U$$1348/X U$$1481/X U$$1614/X VGND VGND VPWR VPWR dadda_fa_1_73_7/CIN
+ dadda_fa_1_72_8/CIN sky130_fd_sc_hd__fa_1
XTAP_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_65_1 U$$536/X U$$669/X U$$802/X VGND VGND VPWR VPWR dadda_fa_1_66_5/CIN
+ dadda_fa_1_65_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_92_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_42_0 dadda_fa_3_42_0/A dadda_fa_3_42_0/B dadda_fa_3_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_0/B dadda_fa_4_42_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_58_0 U$$123/X U$$256/X U$$389/X VGND VGND VPWR VPWR dadda_fa_1_59_6/CIN
+ dadda_fa_1_58_8/A sky130_fd_sc_hd__fa_1
XTAP_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$590 final_adder.U$$598/B final_adder.U$$590/B VGND VGND VPWR VPWR
+ final_adder.U$$710/B sky130_fd_sc_hd__and2_1
XTAP_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$440 U$$440/A U$$474/B VGND VGND VPWR VPWR U$$440/X sky130_fd_sc_hd__xor2_1
XTAP_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$451 U$$40/A1 U$$473/A2 U$$42/A1 U$$473/B2 VGND VGND VPWR VPWR U$$452/A sky130_fd_sc_hd__a22o_1
XTAP_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$462 U$$462/A U$$492/B VGND VGND VPWR VPWR U$$462/X sky130_fd_sc_hd__xor2_1
XFILLER_44_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$473 U$$882/B1 U$$473/A2 U$$64/A1 U$$473/B2 VGND VGND VPWR VPWR U$$474/A sky130_fd_sc_hd__a22o_1
XFILLER_32_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$484 U$$484/A U$$484/B VGND VGND VPWR VPWR U$$484/X sky130_fd_sc_hd__xor2_1
XFILLER_72_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$495 U$$630/B1 U$$537/A2 U$$86/A1 U$$537/B2 VGND VGND VPWR VPWR U$$496/A sky130_fd_sc_hd__a22o_1
XFILLER_72_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_94_3 U$$3919/X U$$4052/X U$$4185/X VGND VGND VPWR VPWR dadda_fa_3_95_1/B
+ dadda_fa_3_94_3/B sky130_fd_sc_hd__fa_1
XFILLER_154_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1340 U$$2797/B VGND VGND VPWR VPWR U$$2755/B sky130_fd_sc_hd__buf_6
XFILLER_160_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1351 U$$184/B VGND VGND VPWR VPWR U$$176/B sky130_fd_sc_hd__buf_4
Xrepeater1362 U$$2716/B VGND VGND VPWR VPWR U$$2739/A sky130_fd_sc_hd__buf_6
Xdadda_fa_2_87_2 U$$4437/X input242/X dadda_fa_2_87_2/CIN VGND VGND VPWR VPWR dadda_fa_3_88_1/A
+ dadda_fa_3_87_3/A sky130_fd_sc_hd__fa_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1373 input31/X VGND VGND VPWR VPWR U$$2569/B sky130_fd_sc_hd__buf_6
XFILLER_99_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1384 U$$2366/B VGND VGND VPWR VPWR U$$2360/B sky130_fd_sc_hd__buf_4
Xdadda_fa_5_64_1 dadda_fa_5_64_1/A dadda_fa_5_64_1/B dadda_fa_5_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_65_0/B dadda_fa_7_64_0/A sky130_fd_sc_hd__fa_2
XFILLER_125_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1395 U$$2303/B VGND VGND VPWR VPWR U$$2273/B sky130_fd_sc_hd__buf_8
XFILLER_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_57_0 dadda_fa_5_57_0/A dadda_fa_5_57_0/B dadda_fa_5_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_58_0/A dadda_fa_6_57_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_56_8 dadda_fa_1_56_8/A dadda_fa_1_56_8/B dadda_fa_1_56_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_57_3/A dadda_fa_3_56_0/A sky130_fd_sc_hd__fa_2
XFILLER_67_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_103_0 U$$2739/Y U$$2873/X U$$3006/X VGND VGND VPWR VPWR dadda_fa_3_104_2/B
+ dadda_fa_3_103_3/B sky130_fd_sc_hd__fa_1
XFILLER_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1190 U$$916/A1 U$$1190/A2 U$$96/A1 U$$1190/B2 VGND VGND VPWR VPWR U$$1191/A sky130_fd_sc_hd__a22o_1
XFILLER_206_1072 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_274 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_82_1 U$$1634/X U$$1767/X U$$1900/X VGND VGND VPWR VPWR dadda_fa_2_83_1/CIN
+ dadda_fa_2_82_4/A sky130_fd_sc_hd__fa_1
XFILLER_85_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_75_0 U$$1620/X U$$1753/X U$$1886/X VGND VGND VPWR VPWR dadda_fa_2_76_0/B
+ dadda_fa_2_75_3/B sky130_fd_sc_hd__fa_1
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_615 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3509 U$$3644/B1 U$$3429/X U$$3511/A1 U$$3430/X VGND VGND VPWR VPWR U$$3510/A sky130_fd_sc_hd__a22o_1
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2808 U$$3356/A1 U$$2810/A2 U$$2808/B1 U$$2810/B2 VGND VGND VPWR VPWR U$$2809/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2819 U$$2819/A U$$2859/B VGND VGND VPWR VPWR U$$2819/X sky130_fd_sc_hd__xor2_1
XFILLER_74_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_102 _346_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 U$$930/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 U$$1746/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 U$$1746/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_422_ _422_/CLK _422_/D VGND VGND VPWR VPWR _422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_179 _197_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_394 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_353_ _355_/CLK _353_/D VGND VGND VPWR VPWR _353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_528 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_284_ _414_/CLK _284_/D VGND VGND VPWR VPWR _284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_97_1 dadda_fa_3_97_1/A dadda_fa_3_97_1/B dadda_fa_3_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_0/CIN dadda_fa_4_97_2/A sky130_fd_sc_hd__fa_1
XFILLER_142_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_74_0 dadda_fa_6_74_0/A dadda_fa_6_74_0/B dadda_fa_6_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_75_0/B dadda_fa_7_74_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_672 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 a[16] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_119_0 U$$3835/Y U$$3969/X U$$4102/X VGND VGND VPWR VPWR dadda_fa_5_120_0/CIN
+ dadda_fa_5_119_1/B sky130_fd_sc_hd__fa_1
XTAP_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$270 U$$270/A U$$272/B VGND VGND VPWR VPWR U$$270/X sky130_fd_sc_hd__xor2_1
XU$$281 U$$281/A U$$317/B VGND VGND VPWR VPWR U$$281/X sky130_fd_sc_hd__xor2_1
XU$$292 U$$703/A1 U$$302/A2 U$$20/A1 U$$302/B2 VGND VGND VPWR VPWR U$$293/A sky130_fd_sc_hd__a22o_1
XFILLER_32_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$6 _302_/Q _174_/Q VGND VGND VPWR VPWR final_adder.U$$6/COUT final_adder.U$$6/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_69_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput301 output301/A VGND VGND VPWR VPWR o[24] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_0 U$$2984/X U$$3117/X U$$3250/X VGND VGND VPWR VPWR dadda_fa_3_93_0/B
+ dadda_fa_3_92_2/B sky130_fd_sc_hd__fa_1
XFILLER_145_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput312 output312/A VGND VGND VPWR VPWR o[34] sky130_fd_sc_hd__buf_2
Xoutput323 output323/A VGND VGND VPWR VPWR o[44] sky130_fd_sc_hd__buf_2
XFILLER_145_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput334 output334/A VGND VGND VPWR VPWR o[54] sky130_fd_sc_hd__buf_2
Xoutput345 output345/A VGND VGND VPWR VPWR o[64] sky130_fd_sc_hd__buf_2
XFILLER_126_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput356 output356/A VGND VGND VPWR VPWR o[74] sky130_fd_sc_hd__buf_2
Xrepeater1170 U$$4418/A1 VGND VGND VPWR VPWR U$$32/B1 sky130_fd_sc_hd__buf_6
Xoutput367 output367/A VGND VGND VPWR VPWR o[84] sky130_fd_sc_hd__buf_2
Xrepeater1181 U$$578/A1 VGND VGND VPWR VPWR U$$850/B1 sky130_fd_sc_hd__buf_6
Xoutput378 output378/A VGND VGND VPWR VPWR o[94] sky130_fd_sc_hd__buf_2
Xdadda_ha_4_118_2 U$$4499/X input149/X VGND VGND VPWR VPWR dadda_fa_5_119_1/A dadda_ha_4_118_2/SUM
+ sky130_fd_sc_hd__ha_1
Xrepeater1192 U$$4410/B1 VGND VGND VPWR VPWR U$$3453/A1 sky130_fd_sc_hd__buf_6
XFILLER_113_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_61_6 dadda_fa_1_61_6/A dadda_fa_1_61_6/B dadda_fa_1_61_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_2/B dadda_fa_2_61_5/B sky130_fd_sc_hd__fa_1
XFILLER_210_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1090 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_5 U$$2775/X U$$2908/X U$$3041/X VGND VGND VPWR VPWR dadda_fa_2_55_2/A
+ dadda_fa_2_54_5/A sky130_fd_sc_hd__fa_1
XFILLER_110_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_47_4 U$$1697/X U$$1830/X U$$1963/X VGND VGND VPWR VPWR dadda_fa_2_48_2/CIN
+ dadda_fa_2_47_5/B sky130_fd_sc_hd__fa_1
XFILLER_167_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_17_2 dadda_fa_4_17_2/A dadda_fa_4_17_2/B dadda_ha_3_17_1/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_18_0/CIN dadda_fa_5_17_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_70_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1020 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_91_0 dadda_fa_7_91_0/A dadda_fa_7_91_0/B dadda_fa_7_91_0/CIN VGND VGND
+ VPWR VPWR _388_/D _259_/D sky130_fd_sc_hd__fa_1
XFILLER_167_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_984 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4007 U$$4418/A1 U$$4043/A2 U$$4420/A1 U$$4043/B2 VGND VGND VPWR VPWR U$$4008/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4018 U$$4018/A U$$4100/B VGND VGND VPWR VPWR U$$4018/X sky130_fd_sc_hd__xor2_1
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4029 U$$4029/A1 U$$4035/A2 U$$4442/A1 U$$4035/B2 VGND VGND VPWR VPWR U$$4030/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3306 U$$3578/B1 U$$3394/A2 U$$431/A1 U$$3394/B2 VGND VGND VPWR VPWR U$$3307/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3317 U$$3317/A U$$3321/B VGND VGND VPWR VPWR U$$3317/X sky130_fd_sc_hd__xor2_1
XFILLER_150_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3328 U$$3737/B1 U$$3348/A2 U$$3876/B1 U$$3346/B2 VGND VGND VPWR VPWR U$$3329/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3339 U$$3339/A U$$3377/B VGND VGND VPWR VPWR U$$3339/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2605 input33/X VGND VGND VPWR VPWR U$$2605/Y sky130_fd_sc_hd__inv_1
XU$$2616 U$$2616/A U$$2624/B VGND VGND VPWR VPWR U$$2616/X sky130_fd_sc_hd__xor2_1
XU$$2627 U$$4269/B1 U$$2683/A2 U$$4408/B1 U$$2683/B2 VGND VGND VPWR VPWR U$$2628/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2638 U$$2638/A U$$2650/B VGND VGND VPWR VPWR U$$2638/X sky130_fd_sc_hd__xor2_1
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1904 U$$1904/A U$$1912/B VGND VGND VPWR VPWR U$$1904/X sky130_fd_sc_hd__xor2_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2649 U$$3880/B1 U$$2653/A2 U$$3747/A1 U$$2653/B2 VGND VGND VPWR VPWR U$$2650/A
+ sky130_fd_sc_hd__a22o_1
XU$$1915 U$$4242/B1 U$$1915/A2 U$$1915/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1916/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1926 U$$2198/B1 U$$1960/A2 U$$2063/B1 U$$1960/B2 VGND VGND VPWR VPWR U$$1927/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1937 U$$1937/A U$$1971/B VGND VGND VPWR VPWR U$$1937/X sky130_fd_sc_hd__xor2_1
XU$$1948 U$$2357/B1 U$$1960/A2 U$$3594/A1 U$$1960/B2 VGND VGND VPWR VPWR U$$1949/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_405_ _407_/CLK _405_/D VGND VGND VPWR VPWR _405_/Q sky130_fd_sc_hd__dfxtp_1
XU$$1959 U$$1959/A U$$2009/B VGND VGND VPWR VPWR U$$1959/X sky130_fd_sc_hd__xor2_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_634 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_336_ _342_/CLK _336_/D VGND VGND VPWR VPWR _336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_267_ _399_/CLK _267_/D VGND VGND VPWR VPWR _267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1019 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_198_ _337_/CLK _198_/D VGND VGND VPWR VPWR _198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_71_5 dadda_fa_2_71_5/A dadda_fa_2_71_5/B dadda_fa_2_71_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_72_2/A dadda_fa_4_71_0/A sky130_fd_sc_hd__fa_1
XFILLER_111_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_634 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_64_4 dadda_fa_2_64_4/A dadda_fa_2_64_4/B dadda_fa_2_64_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_1/CIN dadda_fa_3_64_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater804 U$$2449/B2 VGND VGND VPWR VPWR U$$2459/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater815 U$$2169/B2 VGND VGND VPWR VPWR U$$2091/B2 sky130_fd_sc_hd__buf_4
XFILLER_56_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater826 U$$2046/B2 VGND VGND VPWR VPWR U$$2022/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_57_3 dadda_fa_2_57_3/A dadda_fa_2_57_3/B dadda_fa_2_57_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/B dadda_fa_3_57_3/B sky130_fd_sc_hd__fa_1
Xrepeater837 U$$1869/B2 VGND VGND VPWR VPWR U$$1819/B2 sky130_fd_sc_hd__buf_4
XFILLER_42_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater848 U$$1635/B2 VGND VGND VPWR VPWR U$$1621/B2 sky130_fd_sc_hd__buf_4
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_581 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$11 U$$11/A U$$9/B VGND VGND VPWR VPWR U$$11/X sky130_fd_sc_hd__xor2_1
XFILLER_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater859 U$$259/B2 VGND VGND VPWR VPWR U$$243/B2 sky130_fd_sc_hd__buf_4
XU$$22 U$$22/A1 U$$8/A2 U$$24/A1 U$$8/B2 VGND VGND VPWR VPWR U$$23/A sky130_fd_sc_hd__a22o_1
XU$$33 U$$33/A U$$51/B VGND VGND VPWR VPWR U$$33/X sky130_fd_sc_hd__xor2_1
XU$$44 U$$44/A1 U$$50/A2 U$$44/B1 U$$50/B2 VGND VGND VPWR VPWR U$$45/A sky130_fd_sc_hd__a22o_1
XFILLER_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_27_1 dadda_fa_5_27_1/A dadda_fa_5_27_1/B dadda_fa_5_27_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_28_0/B dadda_fa_7_27_0/A sky130_fd_sc_hd__fa_2
XU$$55 U$$55/A U$$85/B VGND VGND VPWR VPWR U$$55/X sky130_fd_sc_hd__xor2_1
XU$$3840 U$$3838/Y input52/X input51/X U$$3839/X U$$3836/Y VGND VGND VPWR VPWR U$$3840/X
+ sky130_fd_sc_hd__a32o_4
XU$$66 U$$66/A1 U$$98/A2 U$$68/A1 U$$98/B2 VGND VGND VPWR VPWR U$$67/A sky130_fd_sc_hd__a22o_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3851 U$$3851/A U$$3879/B VGND VGND VPWR VPWR U$$3851/X sky130_fd_sc_hd__xor2_1
XFILLER_25_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3862 U$$4273/A1 U$$3902/A2 U$$4273/B1 U$$3902/B2 VGND VGND VPWR VPWR U$$3863/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3873 U$$3873/A U$$3875/B VGND VGND VPWR VPWR U$$3873/X sky130_fd_sc_hd__xor2_1
XU$$77 U$$77/A U$$81/B VGND VGND VPWR VPWR U$$77/X sky130_fd_sc_hd__xor2_1
XFILLER_92_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$88 U$$88/A1 U$$94/A2 U$$90/A1 U$$94/B2 VGND VGND VPWR VPWR U$$89/A sky130_fd_sc_hd__a22o_1
XFILLER_46_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$99 U$$99/A U$$99/B VGND VGND VPWR VPWR U$$99/X sky130_fd_sc_hd__xor2_1
XU$$3884 U$$4293/B1 U$$3970/A2 U$$3884/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3885/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3895 U$$3895/A U$$3909/B VGND VGND VPWR VPWR U$$3895/X sky130_fd_sc_hd__xor2_1
XFILLER_75_1031 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_13 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 _337_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_35 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 _342_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_79 _343_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_101_1 dadda_fa_5_101_1/A dadda_fa_5_101_1/B dadda_fa_5_101_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_102_0/B dadda_fa_7_101_0/A sky130_fd_sc_hd__fa_1
XFILLER_146_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_439 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_39_2 U$$883/X U$$1016/X VGND VGND VPWR VPWR dadda_fa_2_40_4/CIN dadda_fa_3_39_0/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_1_52_2 U$$1175/X U$$1308/X U$$1441/X VGND VGND VPWR VPWR dadda_fa_2_53_1/A
+ dadda_fa_2_52_4/A sky130_fd_sc_hd__fa_1
XFILLER_210_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_45_1 U$$496/X U$$629/X U$$762/X VGND VGND VPWR VPWR dadda_fa_2_46_2/B
+ dadda_fa_2_45_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_22_0 dadda_fa_4_22_0/A dadda_fa_4_22_0/B dadda_fa_4_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/A dadda_fa_5_22_1/A sky130_fd_sc_hd__fa_1
XFILLER_28_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_38_0 U$$83/X U$$216/X U$$349/X VGND VGND VPWR VPWR dadda_fa_2_39_4/B dadda_fa_2_38_5/B
+ sky130_fd_sc_hd__fa_1
XFILLER_102_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1005 final_adder.U$$234/A final_adder.U$$735/X final_adder.U$$235/A2
+ VGND VGND VPWR VPWR final_adder.U$$1045/B sky130_fd_sc_hd__a21o_1
XFILLER_183_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1027 final_adder.U$$3/SUM final_adder.U$$1027/B VGND VGND VPWR VPWR
+ output318/A sky130_fd_sc_hd__xor2_1
XFILLER_137_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$1038 final_adder.U$$240/A final_adder.U$$621/X VGND VGND VPWR VPWR
+ output290/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1049 final_adder.U$$230/B final_adder.U$$1049/B VGND VGND VPWR VPWR
+ output302/A sky130_fd_sc_hd__xor2_1
XFILLER_183_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_670 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_74_3 dadda_fa_3_74_3/A dadda_fa_3_74_3/B dadda_fa_3_74_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_75_1/B dadda_fa_4_74_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_67_2 dadda_fa_3_67_2/A dadda_fa_3_67_2/B dadda_fa_3_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_1/A dadda_fa_4_67_2/B sky130_fd_sc_hd__fa_1
XFILLER_61_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_37_0 dadda_fa_6_37_0/A dadda_fa_6_37_0/B dadda_fa_6_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_38_0/B dadda_fa_7_37_0/CIN sky130_fd_sc_hd__fa_1
XU$$3103 U$$3103/A U$$3109/B VGND VGND VPWR VPWR U$$3103/X sky130_fd_sc_hd__xor2_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3114 U$$3114/A1 U$$3118/A2 U$$3116/A1 U$$3118/B2 VGND VGND VPWR VPWR U$$3115/A
+ sky130_fd_sc_hd__a22o_1
XU$$3125 U$$3125/A U$$3125/B VGND VGND VPWR VPWR U$$3125/X sky130_fd_sc_hd__xor2_1
XU$$3136 input117/X U$$3148/A2 U$$3684/B1 U$$3148/B2 VGND VGND VPWR VPWR U$$3137/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3147 U$$3147/A U$$3150/A VGND VGND VPWR VPWR U$$3147/X sky130_fd_sc_hd__xor2_1
XU$$2402 U$$2402/A U$$2442/B VGND VGND VPWR VPWR U$$2402/X sky130_fd_sc_hd__xor2_1
XU$$2413 U$$3646/A1 U$$2435/A2 U$$3235/B1 U$$2435/B2 VGND VGND VPWR VPWR U$$2414/A
+ sky130_fd_sc_hd__a22o_1
XU$$3158 U$$3158/A U$$3208/B VGND VGND VPWR VPWR U$$3158/X sky130_fd_sc_hd__xor2_1
XU$$3169 U$$3578/B1 U$$3263/A2 U$$431/A1 U$$3263/B2 VGND VGND VPWR VPWR U$$3170/A
+ sky130_fd_sc_hd__a22o_1
XU$$2424 U$$2424/A U$$2454/B VGND VGND VPWR VPWR U$$2424/X sky130_fd_sc_hd__xor2_1
XFILLER_46_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2435 U$$2709/A1 U$$2435/A2 U$$2709/B1 U$$2435/B2 VGND VGND VPWR VPWR U$$2436/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2446 U$$2446/A U$$2446/B VGND VGND VPWR VPWR U$$2446/X sky130_fd_sc_hd__xor2_1
XU$$1701 U$$1701/A U$$1707/B VGND VGND VPWR VPWR U$$1701/X sky130_fd_sc_hd__xor2_1
XFILLER_179_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2457 U$$3416/A1 U$$2459/A2 U$$952/A1 U$$2459/B2 VGND VGND VPWR VPWR U$$2458/A
+ sky130_fd_sc_hd__a22o_1
XU$$1712 U$$2123/A1 U$$1750/A2 U$$1714/A1 U$$1750/B2 VGND VGND VPWR VPWR U$$1713/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2468 input31/X VGND VGND VPWR VPWR U$$2468/Y sky130_fd_sc_hd__inv_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1723 U$$1723/A U$$1751/B VGND VGND VPWR VPWR U$$1723/X sky130_fd_sc_hd__xor2_1
XU$$1734 U$$3102/B1 U$$1736/A2 U$$3243/A1 U$$1736/B2 VGND VGND VPWR VPWR U$$1735/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2479 U$$2479/A U$$2525/B VGND VGND VPWR VPWR U$$2479/X sky130_fd_sc_hd__xor2_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1745 U$$1745/A U$$1780/A VGND VGND VPWR VPWR U$$1745/X sky130_fd_sc_hd__xor2_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1756 U$$660/A1 U$$1764/A2 U$$2717/A1 U$$1764/B2 VGND VGND VPWR VPWR U$$1757/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1767 U$$1767/A U$$1780/A VGND VGND VPWR VPWR U$$1767/X sky130_fd_sc_hd__xor2_1
XFILLER_30_610 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1778 U$$4516/B1 U$$1648/X U$$1778/B1 U$$1649/X VGND VGND VPWR VPWR U$$1779/A sky130_fd_sc_hd__a22o_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1789 U$$2198/B1 U$$1819/A2 U$$2063/B1 U$$1819/B2 VGND VGND VPWR VPWR U$$1790/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_319_ _326_/CLK _319_/D VGND VGND VPWR VPWR _319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput11 a[19] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__buf_6
XFILLER_35_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 a[29] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__buf_6
XFILLER_128_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput33 a[39] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__buf_4
XFILLER_174_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput44 a[49] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_1
Xinput55 a[59] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__buf_6
Xinput66 b[10] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__buf_8
Xinput77 b[20] VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__buf_6
XFILLER_128_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput88 b[30] VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__buf_6
XFILLER_192_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput99 b[40] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__buf_6
XFILLER_170_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_62_1 dadda_fa_2_62_1/A dadda_fa_2_62_1/B dadda_fa_2_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_0/CIN dadda_fa_3_62_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater601 U$$1635/A2 VGND VGND VPWR VPWR U$$1621/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$408 final_adder.U$$412/B final_adder.U$$408/B VGND VGND VPWR VPWR
+ final_adder.U$$532/B sky130_fd_sc_hd__and2_1
Xrepeater612 U$$259/A2 VGND VGND VPWR VPWR U$$243/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$419 final_adder.U$$418/B final_adder.U$$297/X final_adder.U$$293/X
+ VGND VGND VPWR VPWR final_adder.U$$419/X sky130_fd_sc_hd__a21o_1
XFILLER_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater623 U$$1374/X VGND VGND VPWR VPWR U$$1504/A2 sky130_fd_sc_hd__buf_8
XFILLER_38_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_55_0 dadda_fa_2_55_0/A dadda_fa_2_55_0/B dadda_fa_2_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_0/B dadda_fa_3_55_2/B sky130_fd_sc_hd__fa_1
Xrepeater634 U$$1190/A2 VGND VGND VPWR VPWR U$$1174/A2 sky130_fd_sc_hd__buf_6
XFILLER_96_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater645 U$$1083/B2 VGND VGND VPWR VPWR U$$1057/B2 sky130_fd_sc_hd__buf_4
XFILLER_96_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater656 U$$793/B2 VGND VGND VPWR VPWR U$$783/B2 sky130_fd_sc_hd__buf_4
Xrepeater667 U$$678/B2 VGND VGND VPWR VPWR U$$636/B2 sky130_fd_sc_hd__buf_6
XU$$4360 U$$4360/A U$$4366/B VGND VGND VPWR VPWR U$$4360/X sky130_fd_sc_hd__xor2_1
Xrepeater678 U$$491/B2 VGND VGND VPWR VPWR U$$483/B2 sky130_fd_sc_hd__buf_6
Xrepeater689 U$$4226/B2 VGND VGND VPWR VPWR U$$4210/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4371 U$$4508/A1 U$$4373/A2 U$$4510/A1 U$$4373/B2 VGND VGND VPWR VPWR U$$4372/A
+ sky130_fd_sc_hd__a22o_1
XU$$4382 U$$4382/A U$$4382/B VGND VGND VPWR VPWR U$$4382/X sky130_fd_sc_hd__xor2_1
XU$$4393 U$$4393/A U$$4393/B VGND VGND VPWR VPWR U$$4393/X sky130_fd_sc_hd__xor2_1
XFILLER_198_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3670 U$$3944/A1 U$$3686/A2 U$$3944/B1 U$$3686/B2 VGND VGND VPWR VPWR U$$3671/A
+ sky130_fd_sc_hd__a22o_1
XU$$3681 U$$3681/A U$$3683/B VGND VGND VPWR VPWR U$$3681/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3692 U$$4240/A1 U$$3696/A2 U$$4379/A1 U$$3696/B2 VGND VGND VPWR VPWR U$$3693/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_9_0 U$$291/X U$$424/X U$$557/X VGND VGND VPWR VPWR dadda_fa_6_10_0/A dadda_fa_6_9_0/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2980 U$$2980/A input38/X VGND VGND VPWR VPWR U$$2980/X sky130_fd_sc_hd__xor2_1
XFILLER_179_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2991 U$$3813/A1 U$$2995/A2 U$$388/B1 U$$2995/B2 VGND VGND VPWR VPWR U$$2992/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_84_2 dadda_fa_4_84_2/A dadda_fa_4_84_2/B dadda_fa_4_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_85_0/CIN dadda_fa_5_84_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_84_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_77_1 dadda_fa_4_77_1/A dadda_fa_4_77_1/B dadda_fa_4_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/B dadda_fa_5_77_1/B sky130_fd_sc_hd__fa_1
XFILLER_164_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_54_0 dadda_fa_7_54_0/A dadda_fa_7_54_0/B dadda_fa_7_54_0/CIN VGND VGND
+ VPWR VPWR _351_/D _222_/D sky130_fd_sc_hd__fa_1
XTAP_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$931 final_adder.U$$160/A final_adder.U$$869/X final_adder.U$$931/B1
+ VGND VGND VPWR VPWR final_adder.U$$931/X sky130_fd_sc_hd__a21o_1
XTAP_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$953 final_adder.U$$182/A final_adder.U$$891/X final_adder.U$$953/B1
+ VGND VGND VPWR VPWR final_adder.U$$953/X sky130_fd_sc_hd__a21o_1
XU$$803 U$$940/A1 U$$805/A2 U$$940/B1 U$$805/B2 VGND VGND VPWR VPWR U$$804/A sky130_fd_sc_hd__a22o_1
XFILLER_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$975 final_adder.U$$204/A final_adder.U$$817/X final_adder.U$$975/B1
+ VGND VGND VPWR VPWR final_adder.U$$975/X sky130_fd_sc_hd__a21o_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$814 U$$814/A U$$821/A VGND VGND VPWR VPWR U$$814/X sky130_fd_sc_hd__xor2_1
XU$$825 U$$959/A U$$825/B VGND VGND VPWR VPWR U$$825/X sky130_fd_sc_hd__and2_1
XFILLER_16_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$997 final_adder.U$$226/A final_adder.U$$727/X final_adder.U$$997/B1
+ VGND VGND VPWR VPWR final_adder.U$$997/X sky130_fd_sc_hd__a21o_1
XU$$836 U$$836/A1 U$$906/A2 U$$975/A1 U$$906/B2 VGND VGND VPWR VPWR U$$837/A sky130_fd_sc_hd__a22o_1
XU$$847 U$$847/A U$$847/B VGND VGND VPWR VPWR U$$847/X sky130_fd_sc_hd__xor2_1
XU$$858 U$$993/B1 U$$892/A2 U$$997/A1 U$$892/B2 VGND VGND VPWR VPWR U$$859/A sky130_fd_sc_hd__a22o_1
XFILLER_113_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1008 U$$1008/A U$$998/B VGND VGND VPWR VPWR U$$1008/X sky130_fd_sc_hd__xor2_1
XFILLER_71_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$869 U$$869/A U$$877/B VGND VGND VPWR VPWR U$$869/X sky130_fd_sc_hd__xor2_1
XU$$1019 U$$60/A1 U$$993/A2 U$$62/A1 U$$993/B2 VGND VGND VPWR VPWR U$$1020/A sky130_fd_sc_hd__a22o_1
XFILLER_43_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1703 U$$2282/A1 VGND VGND VPWR VPWR U$$90/A1 sky130_fd_sc_hd__buf_4
XFILLER_165_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_72_0 dadda_fa_3_72_0/A dadda_fa_3_72_0/B dadda_fa_3_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_0/B dadda_fa_4_72_1/CIN sky130_fd_sc_hd__fa_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2210 U$$2621/A1 U$$2226/A2 U$$2623/A1 U$$2226/B2 VGND VGND VPWR VPWR U$$2211/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_101_0 dadda_fa_4_101_0/A dadda_fa_4_101_0/B dadda_fa_4_101_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/A dadda_fa_5_101_1/A sky130_fd_sc_hd__fa_1
XU$$2221 U$$2221/A U$$2273/B VGND VGND VPWR VPWR U$$2221/X sky130_fd_sc_hd__xor2_1
XFILLER_47_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_34_5 U$$2336/X U$$2366/B input184/X VGND VGND VPWR VPWR dadda_fa_3_35_2/A
+ dadda_fa_4_34_0/A sky130_fd_sc_hd__fa_1
XU$$2232 U$$4011/B1 U$$2252/A2 U$$4289/A1 U$$2252/B2 VGND VGND VPWR VPWR U$$2233/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2243 U$$2243/A U$$2285/B VGND VGND VPWR VPWR U$$2243/X sky130_fd_sc_hd__xor2_1
XU$$2254 U$$2391/A1 U$$2302/A2 U$$3213/B1 U$$2302/B2 VGND VGND VPWR VPWR U$$2255/A
+ sky130_fd_sc_hd__a22o_1
XU$$2265 U$$2265/A U$$2309/B VGND VGND VPWR VPWR U$$2265/X sky130_fd_sc_hd__xor2_1
XU$$1520 U$$1520/A U$$1546/B VGND VGND VPWR VPWR U$$1520/X sky130_fd_sc_hd__xor2_1
XFILLER_62_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2276 U$$3235/A1 U$$2302/A2 U$$2415/A1 U$$2302/B2 VGND VGND VPWR VPWR U$$2277/A
+ sky130_fd_sc_hd__a22o_1
XU$$1531 U$$1666/B1 U$$1545/A2 U$$985/A1 U$$1545/B2 VGND VGND VPWR VPWR U$$1532/A
+ sky130_fd_sc_hd__a22o_1
XU$$2287 U$$2287/A U$$2328/A VGND VGND VPWR VPWR U$$2287/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1542 U$$1542/A U$$1592/B VGND VGND VPWR VPWR U$$1542/X sky130_fd_sc_hd__xor2_1
XU$$1553 U$$594/A1 U$$1557/A2 U$$594/B1 U$$1557/B2 VGND VGND VPWR VPWR U$$1554/A sky130_fd_sc_hd__a22o_1
XFILLER_37_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2298 U$$2981/B1 U$$2196/X U$$2848/A1 U$$2197/X VGND VGND VPWR VPWR U$$2299/A sky130_fd_sc_hd__a22o_1
XU$$1564 U$$1564/A U$$1592/B VGND VGND VPWR VPWR U$$1564/X sky130_fd_sc_hd__xor2_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1575 U$$342/A1 U$$1575/A2 U$$1714/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1576/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1586 U$$1586/A U$$1620/B VGND VGND VPWR VPWR U$$1586/X sky130_fd_sc_hd__xor2_1
XFILLER_124_1113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1597 U$$2282/A1 U$$1607/A2 U$$2967/B1 U$$1607/B2 VGND VGND VPWR VPWR U$$1598/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_94_1 dadda_fa_5_94_1/A dadda_fa_5_94_1/B dadda_fa_5_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_95_0/B dadda_fa_7_94_0/A sky130_fd_sc_hd__fa_1
XFILLER_147_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_87_0 dadda_fa_5_87_0/A dadda_fa_5_87_0/B dadda_fa_5_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_88_0/A dadda_fa_6_87_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_79_7 U$$3889/X U$$4022/X U$$4155/X VGND VGND VPWR VPWR dadda_fa_2_80_2/CIN
+ dadda_fa_2_79_5/CIN sky130_fd_sc_hd__fa_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4433_1793 VGND VGND VPWR VPWR U$$4433_1793/HI U$$4433/B sky130_fd_sc_hd__conb_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$205 final_adder.U$$204/B final_adder.U$$975/B1 final_adder.U$$205/B1
+ VGND VGND VPWR VPWR final_adder.U$$205/X sky130_fd_sc_hd__a21o_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$216 final_adder.U$$216/A final_adder.U$$216/B VGND VGND VPWR VPWR
+ final_adder.U$$344/B sky130_fd_sc_hd__and2_1
Xrepeater420 U$$4369/A2 VGND VGND VPWR VPWR U$$4361/A2 sky130_fd_sc_hd__buf_4
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$227 final_adder.U$$226/B final_adder.U$$997/B1 final_adder.U$$227/B1
+ VGND VGND VPWR VPWR final_adder.U$$227/X sky130_fd_sc_hd__a21o_1
Xrepeater431 U$$4164/A2 VGND VGND VPWR VPWR U$$4144/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$238 final_adder.U$$238/A final_adder.U$$238/B VGND VGND VPWR VPWR
+ final_adder.U$$366/B sky130_fd_sc_hd__and2_1
XTAP_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater442 U$$80/A2 VGND VGND VPWR VPWR U$$50/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$249 final_adder.U$$7/SUM final_adder.U$$6/COUT final_adder.U$$7/COUT
+ VGND VGND VPWR VPWR final_adder.U$$249/X sky130_fd_sc_hd__a21o_1
Xrepeater453 U$$3977/X VGND VGND VPWR VPWR U$$4101/A2 sky130_fd_sc_hd__buf_6
Xrepeater464 U$$3777/A2 VGND VGND VPWR VPWR U$$3753/A2 sky130_fd_sc_hd__buf_6
Xrepeater475 U$$3696/A2 VGND VGND VPWR VPWR U$$3686/A2 sky130_fd_sc_hd__buf_6
XFILLER_27_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater486 U$$3429/X VGND VGND VPWR VPWR U$$3517/A2 sky130_fd_sc_hd__buf_6
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater497 U$$3255/A2 VGND VGND VPWR VPWR U$$3285/A2 sky130_fd_sc_hd__buf_6
XU$$4509_1831 VGND VGND VPWR VPWR U$$4509_1831/HI U$$4509/B sky130_fd_sc_hd__conb_1
XU$$4190 U$$4464/A1 U$$4210/A2 U$$4466/A1 U$$4210/B2 VGND VGND VPWR VPWR U$$4191/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_103_2 dadda_fa_3_103_2/A dadda_fa_3_103_2/B dadda_fa_3_103_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_104_1/A dadda_fa_4_103_2/B sky130_fd_sc_hd__fa_1
XFILLER_88_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput201 c[4] VGND VGND VPWR VPWR input201/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput212 c[5] VGND VGND VPWR VPWR input212/X sky130_fd_sc_hd__buf_4
XFILLER_49_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput223 c[6] VGND VGND VPWR VPWR input223/X sky130_fd_sc_hd__clkbuf_4
XTAP_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput234 c[7] VGND VGND VPWR VPWR input234/X sky130_fd_sc_hd__clkbuf_4
XTAP_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 c[8] VGND VGND VPWR VPWR input245/X sky130_fd_sc_hd__clkbuf_4
XFILLER_48_326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_67_5 U$$2136/X U$$2269/X U$$2402/X VGND VGND VPWR VPWR dadda_fa_1_68_7/A
+ dadda_fa_2_67_0/A sky130_fd_sc_hd__fa_1
Xinput256 c[9] VGND VGND VPWR VPWR input256/X sky130_fd_sc_hd__buf_4
XTAP_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_117_0 dadda_fa_6_117_0/A dadda_fa_6_117_0/B dadda_fa_6_117_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_118_0/B dadda_fa_7_117_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$750 final_adder.U$$782/B final_adder.U$$750/B VGND VGND VPWR VPWR
+ final_adder.U$$750/X sky130_fd_sc_hd__and2_1
XTAP_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$761 final_adder.U$$760/B final_adder.U$$681/X final_adder.U$$649/X
+ VGND VGND VPWR VPWR final_adder.U$$761/X sky130_fd_sc_hd__a21o_1
XTAP_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$600 U$$52/A1 U$$616/A2 U$$52/B1 U$$616/B2 VGND VGND VPWR VPWR U$$601/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$772 final_adder.U$$772/A final_adder.U$$772/B VGND VGND VPWR VPWR
+ final_adder.U$$772/X sky130_fd_sc_hd__and2_1
XTAP_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$611 U$$611/A U$$637/B VGND VGND VPWR VPWR U$$611/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$783 final_adder.U$$782/B final_adder.U$$703/X final_adder.U$$671/X
+ VGND VGND VPWR VPWR final_adder.U$$783/X sky130_fd_sc_hd__a21o_1
XU$$622 U$$896/A1 U$$624/A2 U$$759/B1 U$$624/B2 VGND VGND VPWR VPWR U$$623/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_37_3 dadda_fa_3_37_3/A dadda_fa_3_37_3/B dadda_fa_3_37_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_38_1/B dadda_fa_4_37_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$794 final_adder.U$$794/A final_adder.U$$794/B VGND VGND VPWR VPWR
+ final_adder.U$$794/X sky130_fd_sc_hd__and2_1
XU$$633 U$$633/A U$$637/B VGND VGND VPWR VPWR U$$633/X sky130_fd_sc_hd__xor2_1
XU$$644 U$$918/A1 U$$652/A2 U$$920/A1 U$$652/B2 VGND VGND VPWR VPWR U$$645/A sky130_fd_sc_hd__a22o_1
XFILLER_90_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$655 U$$655/A U$$684/A VGND VGND VPWR VPWR U$$655/X sky130_fd_sc_hd__xor2_1
XU$$666 U$$940/A1 U$$672/A2 U$$940/B1 U$$668/B2 VGND VGND VPWR VPWR U$$667/A sky130_fd_sc_hd__a22o_1
XFILLER_95_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$677 U$$677/A U$$683/B VGND VGND VPWR VPWR U$$677/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$688 input3/X U$$688/B VGND VGND VPWR VPWR U$$688/X sky130_fd_sc_hd__and2_1
XFILLER_182_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$699 U$$836/A1 U$$711/A2 U$$975/A1 U$$711/B2 VGND VGND VPWR VPWR U$$700/A sky130_fd_sc_hd__a22o_1
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1500 U$$4103/B1 VGND VGND VPWR VPWR U$$2324/A1 sky130_fd_sc_hd__buf_4
Xrepeater1511 U$$4240/A1 VGND VGND VPWR VPWR U$$3829/A1 sky130_fd_sc_hd__buf_4
Xrepeater1522 U$$18/A1 VGND VGND VPWR VPWR U$$703/A1 sky130_fd_sc_hd__buf_6
Xrepeater1533 U$$111/B VGND VGND VPWR VPWR U$$81/B sky130_fd_sc_hd__buf_6
XFILLER_181_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1544 input119/X VGND VGND VPWR VPWR U$$3960/B1 sky130_fd_sc_hd__buf_4
Xrepeater1555 U$$3684/A1 VGND VGND VPWR VPWR U$$122/A1 sky130_fd_sc_hd__buf_6
XFILLER_153_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1566 U$$2312/A1 VGND VGND VPWR VPWR U$$940/B1 sky130_fd_sc_hd__buf_4
XFILLER_119_1215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1577 input115/X VGND VGND VPWR VPWR U$$4228/A1 sky130_fd_sc_hd__buf_4
XFILLER_154_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1588 U$$2032/A1 VGND VGND VPWR VPWR U$$799/A1 sky130_fd_sc_hd__buf_6
XFILLER_98_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1599 U$$2715/A1 VGND VGND VPWR VPWR U$$660/A1 sky130_fd_sc_hd__buf_8
XFILLER_98_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_32_2 U$$869/X U$$1002/X U$$1135/X VGND VGND VPWR VPWR dadda_fa_3_33_1/A
+ dadda_fa_3_32_3/A sky130_fd_sc_hd__fa_1
XU$$2040 U$$2312/B1 U$$2040/A2 U$$807/B1 U$$2040/B2 VGND VGND VPWR VPWR U$$2041/A
+ sky130_fd_sc_hd__a22o_1
XU$$2051 U$$2051/A U$$2054/A VGND VGND VPWR VPWR U$$2051/X sky130_fd_sc_hd__xor2_1
XU$$2062 U$$2062/A U$$2094/B VGND VGND VPWR VPWR U$$2062/X sky130_fd_sc_hd__xor2_1
XU$$2073 U$$2621/A1 U$$2099/A2 U$$3719/A1 U$$2099/B2 VGND VGND VPWR VPWR U$$2074/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2084 U$$2084/A U$$2092/B VGND VGND VPWR VPWR U$$2084/X sky130_fd_sc_hd__xor2_1
XFILLER_23_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1350 U$$1350/A U$$1354/B VGND VGND VPWR VPWR U$$1350/X sky130_fd_sc_hd__xor2_1
XU$$2095 U$$4011/B1 U$$2099/A2 U$$864/A1 U$$2099/B2 VGND VGND VPWR VPWR U$$2096/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1361 U$$2318/B1 U$$1361/A2 U$$952/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1362/A
+ sky130_fd_sc_hd__a22o_1
XU$$1372 U$$1506/A VGND VGND VPWR VPWR U$$1372/Y sky130_fd_sc_hd__inv_1
XFILLER_50_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1383 U$$1383/A U$$1405/B VGND VGND VPWR VPWR U$$1383/X sky130_fd_sc_hd__xor2_1
XFILLER_188_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1394 U$$1666/B1 U$$1422/A2 U$$985/A1 U$$1422/B2 VGND VGND VPWR VPWR U$$1395/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_106_0_1863 VGND VGND VPWR VPWR dadda_fa_2_106_0/A dadda_fa_2_106_0_1863/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_108_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_84_5 U$$3367/X U$$3500/X U$$3633/X VGND VGND VPWR VPWR dadda_fa_2_85_3/CIN
+ dadda_fa_2_84_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_77_4 U$$2954/X U$$3087/X U$$3220/X VGND VGND VPWR VPWR dadda_fa_2_78_1/CIN
+ dadda_fa_2_77_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_47_2 dadda_fa_4_47_2/A dadda_fa_4_47_2/B dadda_fa_4_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_48_0/CIN dadda_fa_5_47_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_476 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_17_0 dadda_fa_7_17_0/A dadda_fa_7_17_0/B dadda_fa_7_17_0/CIN VGND VGND
+ VPWR VPWR _314_/D _185_/D sky130_fd_sc_hd__fa_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$90 _386_/Q _258_/Q VGND VGND VPWR VPWR final_adder.U$$935/B1 final_adder.U$$164/A
+ sky130_fd_sc_hd__ha_1
XFILLER_201_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_754 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_894 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_73 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_59_3 U$$1322/X U$$1455/X VGND VGND VPWR VPWR dadda_fa_1_60_7/B dadda_fa_2_59_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_95_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_70_0_1848 VGND VGND VPWR VPWR dadda_fa_0_70_0/A dadda_fa_0_70_0_1848/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_27_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_65_2 U$$935/X U$$1068/X U$$1201/X VGND VGND VPWR VPWR dadda_fa_1_66_6/A
+ dadda_fa_1_65_8/A sky130_fd_sc_hd__fa_1
XTAP_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_42_1 dadda_fa_3_42_1/A dadda_fa_3_42_1/B dadda_fa_3_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_0/CIN dadda_fa_4_42_2/A sky130_fd_sc_hd__fa_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_58_1 U$$522/X U$$655/X U$$788/X VGND VGND VPWR VPWR dadda_fa_1_59_7/A
+ dadda_fa_1_58_8/B sky130_fd_sc_hd__fa_1
XTAP_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$580 final_adder.U$$588/B final_adder.U$$580/B VGND VGND VPWR VPWR
+ final_adder.U$$700/B sky130_fd_sc_hd__and2_1
XTAP_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_35_0 dadda_fa_3_35_0/A dadda_fa_3_35_0/B dadda_fa_3_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_0/B dadda_fa_4_35_1/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$591 final_adder.U$$590/B final_adder.U$$475/X final_adder.U$$467/X
+ VGND VGND VPWR VPWR final_adder.U$$591/X sky130_fd_sc_hd__a21o_1
XU$$430 U$$430/A U$$516/B VGND VGND VPWR VPWR U$$430/X sky130_fd_sc_hd__xor2_1
XTAP_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$441 U$$850/B1 U$$473/A2 U$$717/A1 U$$473/B2 VGND VGND VPWR VPWR U$$442/A sky130_fd_sc_hd__a22o_1
XFILLER_189_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$452 U$$452/A U$$474/B VGND VGND VPWR VPWR U$$452/X sky130_fd_sc_hd__xor2_1
XFILLER_204_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$463 U$$463/A1 U$$483/A2 U$$54/A1 U$$483/B2 VGND VGND VPWR VPWR U$$464/A sky130_fd_sc_hd__a22o_1
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$474 U$$474/A U$$474/B VGND VGND VPWR VPWR U$$474/X sky130_fd_sc_hd__xor2_1
XU$$485 U$$896/A1 U$$491/A2 U$$759/B1 U$$491/B2 VGND VGND VPWR VPWR U$$486/A sky130_fd_sc_hd__a22o_1
XU$$496 U$$496/A U$$536/B VGND VGND VPWR VPWR U$$496/X sky130_fd_sc_hd__xor2_1
XFILLER_32_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_1206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_94_4 U$$4318/X U$$4451/X input250/X VGND VGND VPWR VPWR dadda_fa_3_95_1/CIN
+ dadda_fa_3_94_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1330 input40/X VGND VGND VPWR VPWR U$$3151/A sky130_fd_sc_hd__buf_4
XFILLER_114_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1341 U$$2825/B VGND VGND VPWR VPWR U$$2797/B sky130_fd_sc_hd__buf_6
XFILLER_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1352 U$$212/B VGND VGND VPWR VPWR U$$184/B sky130_fd_sc_hd__buf_4
XFILLER_114_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_87_3 dadda_fa_2_87_3/A dadda_fa_2_87_3/B dadda_fa_2_87_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_1/B dadda_fa_3_87_3/B sky130_fd_sc_hd__fa_1
Xrepeater1363 U$$2710/B VGND VGND VPWR VPWR U$$2680/B sky130_fd_sc_hd__buf_8
Xrepeater1374 input31/X VGND VGND VPWR VPWR U$$2603/A sky130_fd_sc_hd__buf_4
XFILLER_99_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1385 U$$2426/B VGND VGND VPWR VPWR U$$2366/B sky130_fd_sc_hd__buf_8
Xrepeater1396 U$$2328/A VGND VGND VPWR VPWR U$$2285/B sky130_fd_sc_hd__buf_6
XFILLER_140_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_57_1 dadda_fa_5_57_1/A dadda_fa_5_57_1/B dadda_fa_5_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_58_0/B dadda_fa_7_57_0/A sky130_fd_sc_hd__fa_2
XFILLER_68_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_103_1 U$$3139/X U$$3272/X U$$3405/X VGND VGND VPWR VPWR dadda_fa_3_104_2/CIN
+ dadda_fa_3_103_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_23_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1180 U$$4055/B1 U$$1222/A2 U$$3922/A1 U$$1222/B2 VGND VGND VPWR VPWR U$$1181/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1191 U$$1191/A U$$1209/B VGND VGND VPWR VPWR U$$1191/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_124_0 dadda_fa_5_124_0/A U$$4245/X U$$4378/X VGND VGND VPWR VPWR dadda_fa_6_125_0/B
+ dadda_fa_6_124_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_206_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_82_2 U$$2033/X U$$2166/X U$$2299/X VGND VGND VPWR VPWR dadda_fa_2_83_2/A
+ dadda_fa_2_82_4/B sky130_fd_sc_hd__fa_1
XFILLER_78_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1099 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_75_1 U$$2019/X U$$2152/X U$$2285/X VGND VGND VPWR VPWR dadda_fa_2_76_0/CIN
+ dadda_fa_2_75_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_52_0 dadda_fa_4_52_0/A dadda_fa_4_52_0/B dadda_fa_4_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/A dadda_fa_5_52_1/A sky130_fd_sc_hd__fa_1
XFILLER_58_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_68_0 U$$2537/X U$$2670/X U$$2803/X VGND VGND VPWR VPWR dadda_fa_2_69_0/B
+ dadda_fa_2_68_3/B sky130_fd_sc_hd__fa_1
Xdadda_ha_2_102_3 U$$3802/X U$$3935/X VGND VGND VPWR VPWR dadda_fa_3_103_3/A dadda_fa_4_102_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_19_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2809 U$$2809/A U$$2817/B VGND VGND VPWR VPWR U$$2809/X sky130_fd_sc_hd__xor2_1
XFILLER_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _384_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _390_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 U$$930/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_421_ _421_/CLK _421_/D VGND VGND VPWR VPWR _421_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_183_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 U$$217/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_158 U$$98/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_169 _196_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_352_ _355_/CLK _352_/D VGND VGND VPWR VPWR _352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_283_ _412_/CLK _283_/D VGND VGND VPWR VPWR _283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_97_2 dadda_fa_3_97_2/A dadda_fa_3_97_2/B dadda_fa_3_97_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_1/A dadda_fa_4_97_2/B sky130_fd_sc_hd__fa_1
XFILLER_68_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_67_0 dadda_fa_6_67_0/A dadda_fa_6_67_0/B dadda_fa_6_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_68_0/B dadda_fa_7_67_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_146_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_70_0 dadda_fa_0_70_0/A U$$546/X U$$679/X VGND VGND VPWR VPWR dadda_fa_1_71_6/B
+ dadda_fa_1_70_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 a[17] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_4
XTAP_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_119_1 U$$4235/X U$$4368/X U$$4501/X VGND VGND VPWR VPWR dadda_fa_5_120_1/A
+ dadda_fa_5_119_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_5_6_1 U$$418/X U$$436/B VGND VGND VPWR VPWR dadda_fa_6_7_0/B dadda_fa_7_6_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$260 U$$260/A U$$260/B VGND VGND VPWR VPWR U$$260/X sky130_fd_sc_hd__xor2_1
XFILLER_91_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$271 U$$817/B1 U$$141/X U$$271/B1 U$$142/X VGND VGND VPWR VPWR U$$272/A sky130_fd_sc_hd__a22o_1
XFILLER_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$282 U$$8/A1 U$$316/A2 U$$8/B1 U$$316/B2 VGND VGND VPWR VPWR U$$283/A sky130_fd_sc_hd__a22o_1
XU$$293 U$$293/A U$$379/B VGND VGND VPWR VPWR U$$293/X sky130_fd_sc_hd__xor2_1
XFILLER_162_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_691 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$7 _303_/Q _175_/Q VGND VGND VPWR VPWR final_adder.U$$7/COUT final_adder.U$$7/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_195_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput302 output302/A VGND VGND VPWR VPWR o[25] sky130_fd_sc_hd__buf_2
XFILLER_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_92_1 U$$3383/X U$$3516/X U$$3649/X VGND VGND VPWR VPWR dadda_fa_3_93_0/CIN
+ dadda_fa_3_92_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_127_982 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput313 output313/A VGND VGND VPWR VPWR o[35] sky130_fd_sc_hd__buf_2
XFILLER_133_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput324 output324/A VGND VGND VPWR VPWR o[45] sky130_fd_sc_hd__buf_2
Xoutput335 output335/A VGND VGND VPWR VPWR o[55] sky130_fd_sc_hd__buf_2
Xoutput346 output346/A VGND VGND VPWR VPWR o[65] sky130_fd_sc_hd__buf_2
XFILLER_160_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1160 U$$1076/B VGND VGND VPWR VPWR U$$1095/A sky130_fd_sc_hd__buf_8
Xdadda_fa_2_85_0 U$$3901/X U$$4034/X U$$4167/X VGND VGND VPWR VPWR dadda_fa_3_86_0/B
+ dadda_fa_3_85_2/B sky130_fd_sc_hd__fa_1
XFILLER_114_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1171 input69/X VGND VGND VPWR VPWR U$$4418/A1 sky130_fd_sc_hd__buf_4
XFILLER_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput357 output357/A VGND VGND VPWR VPWR o[75] sky130_fd_sc_hd__buf_2
XFILLER_160_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput368 output368/A VGND VGND VPWR VPWR o[85] sky130_fd_sc_hd__buf_2
Xrepeater1182 U$$578/A1 VGND VGND VPWR VPWR U$$989/A1 sky130_fd_sc_hd__buf_8
Xoutput379 output379/A VGND VGND VPWR VPWR o[95] sky130_fd_sc_hd__buf_2
Xrepeater1193 U$$4410/B1 VGND VGND VPWR VPWR U$$711/B1 sky130_fd_sc_hd__buf_6
XFILLER_206_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_48_7 U$$2896/X U$$3029/X VGND VGND VPWR VPWR dadda_fa_2_49_3/B dadda_fa_3_48_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_102_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_7 dadda_fa_1_61_7/A dadda_fa_1_61_7/B dadda_fa_1_61_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_2/CIN dadda_fa_2_61_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_171_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_6 U$$3174/X U$$3307/X U$$3440/X VGND VGND VPWR VPWR dadda_fa_2_55_2/B
+ dadda_fa_2_54_5/B sky130_fd_sc_hd__fa_1
XFILLER_132_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_958 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_47_5 U$$2096/X U$$2229/X U$$2362/X VGND VGND VPWR VPWR dadda_fa_2_48_3/A
+ dadda_fa_2_47_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_167_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_6_0 dadda_fa_7_6_0/A dadda_fa_7_6_0/B dadda_fa_7_6_0/CIN VGND VGND VPWR
+ VPWR _303_/D _174_/D sky130_fd_sc_hd__fa_1
XFILLER_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_595 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_84_0 dadda_fa_7_84_0/A dadda_fa_7_84_0/B dadda_fa_7_84_0/CIN VGND VGND
+ VPWR VPWR _381_/D _252_/D sky130_fd_sc_hd__fa_2
XFILLER_178_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4008 U$$4008/A U$$4044/B VGND VGND VPWR VPWR U$$4008/X sky130_fd_sc_hd__xor2_1
XU$$4019 U$$4019/A1 U$$4107/A2 U$$4293/B1 U$$4107/B2 VGND VGND VPWR VPWR U$$4020/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3307 U$$3307/A U$$3395/B VGND VGND VPWR VPWR U$$3307/X sky130_fd_sc_hd__xor2_1
XFILLER_19_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3318 U$$989/A1 U$$3320/A2 U$$991/A1 U$$3320/B2 VGND VGND VPWR VPWR U$$3319/A sky130_fd_sc_hd__a22o_1
XU$$3329 U$$3329/A U$$3349/B VGND VGND VPWR VPWR U$$3329/X sky130_fd_sc_hd__xor2_1
XFILLER_18_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2606 input33/X U$$2606/B VGND VGND VPWR VPWR U$$2606/X sky130_fd_sc_hd__and2_1
XU$$2617 U$$3028/A1 U$$2625/A2 U$$2754/B1 U$$2625/B2 VGND VGND VPWR VPWR U$$2618/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2628 U$$2628/A U$$2658/B VGND VGND VPWR VPWR U$$2628/X sky130_fd_sc_hd__xor2_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2639 U$$4146/A1 U$$2727/A2 input71/X U$$2727/B2 VGND VGND VPWR VPWR U$$2640/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1905 U$$807/B1 U$$1785/X U$$948/A1 U$$1786/X VGND VGND VPWR VPWR U$$1906/A sky130_fd_sc_hd__a22o_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1916 U$$1916/A U$$1917/A VGND VGND VPWR VPWR U$$1916/X sky130_fd_sc_hd__xor2_1
XFILLER_33_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1927 U$$1927/A U$$1993/B VGND VGND VPWR VPWR U$$1927/X sky130_fd_sc_hd__xor2_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clkbuf_3_1_0_clk/X VGND VGND VPWR VPWR _360_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1938 U$$4404/A1 U$$1970/A2 U$$981/A1 U$$1970/B2 VGND VGND VPWR VPWR U$$1939/A
+ sky130_fd_sc_hd__a22o_1
X_404_ _407_/CLK _404_/D VGND VGND VPWR VPWR _404_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1949 U$$1949/A U$$1993/B VGND VGND VPWR VPWR U$$1949/X sky130_fd_sc_hd__xor2_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_335_ _337_/CLK _335_/D VGND VGND VPWR VPWR _335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_266_ _399_/CLK _266_/D VGND VGND VPWR VPWR _266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_197_ _329_/CLK _197_/D VGND VGND VPWR VPWR _197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_64_5 dadda_fa_2_64_5/A dadda_fa_2_64_5/B dadda_fa_2_64_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_65_2/A dadda_fa_4_64_0/A sky130_fd_sc_hd__fa_2
XFILLER_111_646 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater805 U$$2334/X VGND VGND VPWR VPWR U$$2449/B2 sky130_fd_sc_hd__buf_6
Xrepeater816 U$$2099/B2 VGND VGND VPWR VPWR U$$2113/B2 sky130_fd_sc_hd__buf_4
XFILLER_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater827 U$$2046/B2 VGND VGND VPWR VPWR U$$2052/B2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_57_4 dadda_fa_2_57_4/A dadda_fa_2_57_4/B dadda_fa_2_57_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_1/CIN dadda_fa_3_57_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater838 U$$1786/X VGND VGND VPWR VPWR U$$1869/B2 sky130_fd_sc_hd__clkbuf_8
Xrepeater849 U$$1637/B2 VGND VGND VPWR VPWR U$$1635/B2 sky130_fd_sc_hd__buf_6
XU$$12 U$$12/A1 U$$8/A2 U$$14/A1 U$$8/B2 VGND VGND VPWR VPWR U$$13/A sky130_fd_sc_hd__a22o_1
XFILLER_77_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$23 U$$23/A U$$9/B VGND VGND VPWR VPWR U$$23/X sky130_fd_sc_hd__xor2_1
XFILLER_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$34 U$$34/A1 U$$50/A2 U$$36/A1 U$$50/B2 VGND VGND VPWR VPWR U$$35/A sky130_fd_sc_hd__a22o_1
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3830 U$$3830/A U$$3834/B VGND VGND VPWR VPWR U$$3830/X sky130_fd_sc_hd__xor2_1
XU$$45 U$$45/A U$$51/B VGND VGND VPWR VPWR U$$45/X sky130_fd_sc_hd__xor2_1
XU$$3841 U$$3839/B input51/X input52/X U$$3836/Y VGND VGND VPWR VPWR U$$3841/X sky130_fd_sc_hd__a22o_4
XTAP_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$56 U$$56/A1 U$$98/A2 U$$56/B1 U$$98/B2 VGND VGND VPWR VPWR U$$57/A sky130_fd_sc_hd__a22o_1
XU$$3852 U$$3852/A1 U$$3874/A2 U$$3852/B1 U$$3874/B2 VGND VGND VPWR VPWR U$$3853/A
+ sky130_fd_sc_hd__a22o_1
XU$$67 U$$67/A U$$85/B VGND VGND VPWR VPWR U$$67/X sky130_fd_sc_hd__xor2_1
XU$$3863 U$$3863/A U$$3903/B VGND VGND VPWR VPWR U$$3863/X sky130_fd_sc_hd__xor2_1
XU$$78 U$$78/A1 U$$80/A2 U$$80/A1 U$$80/B2 VGND VGND VPWR VPWR U$$79/A sky130_fd_sc_hd__a22o_1
XU$$3874 U$$4422/A1 U$$3874/A2 U$$4424/A1 U$$3874/B2 VGND VGND VPWR VPWR U$$3875/A
+ sky130_fd_sc_hd__a22o_1
XU$$89 U$$89/A U$$99/B VGND VGND VPWR VPWR U$$89/X sky130_fd_sc_hd__xor2_1
XFILLER_64_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3885 U$$3885/A U$$3971/B VGND VGND VPWR VPWR U$$3885/X sky130_fd_sc_hd__xor2_1
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3896 U$$4442/B1 U$$3902/A2 U$$4309/A1 U$$3902/B2 VGND VGND VPWR VPWR U$$3897/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_clk _385_/CLK VGND VGND VPWR VPWR _423_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1043 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1002 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1087 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_14 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 _337_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_36 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_69 _342_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_52_3 U$$1574/X U$$1707/X U$$1840/X VGND VGND VPWR VPWR dadda_fa_2_53_1/B
+ dadda_fa_2_52_4/B sky130_fd_sc_hd__fa_1
XFILLER_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_45_2 U$$895/X U$$1028/X U$$1161/X VGND VGND VPWR VPWR dadda_fa_2_46_2/CIN
+ dadda_fa_2_45_5/A sky130_fd_sc_hd__fa_1
XFILLER_16_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_22_1 dadda_fa_4_22_1/A dadda_fa_4_22_1/B dadda_fa_4_22_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/B dadda_fa_5_22_1/B sky130_fd_sc_hd__fa_1
XFILLER_83_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_38_1 U$$482/X U$$615/X U$$748/X VGND VGND VPWR VPWR dadda_fa_2_39_4/CIN
+ dadda_fa_2_38_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_110_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_clk _380_/CLK VGND VGND VPWR VPWR _381_/CLK sky130_fd_sc_hd__clkbuf_16
Xdadda_fa_4_15_0 U$$303/X U$$436/X U$$569/X VGND VGND VPWR VPWR dadda_fa_5_16_0/A
+ dadda_fa_5_15_1/A sky130_fd_sc_hd__fa_1
XFILLER_52_950 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1017 final_adder.U$$8/SUM final_adder.U$$503/X final_adder.U$$8/COUT
+ VGND VGND VPWR VPWR final_adder.U$$1033/B sky130_fd_sc_hd__a21o_1
XFILLER_183_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1028 final_adder.U$$4/SUM final_adder.U$$381/X VGND VGND VPWR VPWR
+ output329/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1039 final_adder.U$$240/B final_adder.U$$1039/B VGND VGND VPWR VPWR
+ output291/A sky130_fd_sc_hd__xor2_1
XFILLER_165_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_833 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_67_3 dadda_fa_3_67_3/A dadda_fa_3_67_3/B dadda_fa_3_67_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_68_1/B dadda_fa_4_67_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_87_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3104 U$$3378/A1 U$$3108/A2 U$$3243/A1 U$$3108/B2 VGND VGND VPWR VPWR U$$3105/A
+ sky130_fd_sc_hd__a22o_1
XU$$3115 U$$3115/A U$$3117/B VGND VGND VPWR VPWR U$$3115/X sky130_fd_sc_hd__xor2_1
XU$$3126 U$$384/B1 U$$3132/A2 U$$251/A1 U$$3132/B2 VGND VGND VPWR VPWR U$$3127/A sky130_fd_sc_hd__a22o_1
XFILLER_19_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3137 U$$3137/A U$$3150/A VGND VGND VPWR VPWR U$$3137/X sky130_fd_sc_hd__xor2_1
XFILLER_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3148 U$$3148/A1 U$$3148/A2 U$$3148/B1 U$$3148/B2 VGND VGND VPWR VPWR U$$3149/A
+ sky130_fd_sc_hd__a22o_1
XU$$2403 U$$3499/A1 U$$2403/A2 U$$896/B1 U$$2403/B2 VGND VGND VPWR VPWR U$$2404/A
+ sky130_fd_sc_hd__a22o_1
XU$$3159 U$$3159/A1 U$$3207/A2 U$$3159/B1 U$$3207/B2 VGND VGND VPWR VPWR U$$3160/A
+ sky130_fd_sc_hd__a22o_1
XU$$2414 U$$2414/A U$$2446/B VGND VGND VPWR VPWR U$$2414/X sky130_fd_sc_hd__xor2_1
XFILLER_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2425 U$$2425/A1 U$$2435/A2 U$$4480/B1 U$$2435/B2 VGND VGND VPWR VPWR U$$2426/A
+ sky130_fd_sc_hd__a22o_1
XU$$2436 U$$2436/A U$$2446/B VGND VGND VPWR VPWR U$$2436/X sky130_fd_sc_hd__xor2_1
XFILLER_36_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1702 U$$878/B1 U$$1706/A2 U$$2113/B1 U$$1706/B2 VGND VGND VPWR VPWR U$$1703/A
+ sky130_fd_sc_hd__a22o_1
XU$$2447 U$$4228/A1 U$$2449/A2 U$$4365/B1 U$$2449/B2 VGND VGND VPWR VPWR U$$2448/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2458 U$$2458/A U$$2465/A VGND VGND VPWR VPWR U$$2458/X sky130_fd_sc_hd__xor2_1
XU$$1713 U$$1713/A U$$1721/B VGND VGND VPWR VPWR U$$1713/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_26_clk _380_/CLK VGND VGND VPWR VPWR _407_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$1724 U$$3366/B1 U$$1736/A2 U$$2409/B1 U$$1736/B2 VGND VGND VPWR VPWR U$$1725/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2469 input31/X U$$2469/B VGND VGND VPWR VPWR U$$2469/X sky130_fd_sc_hd__and2_1
XFILLER_62_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1735 U$$1735/A U$$1779/B VGND VGND VPWR VPWR U$$1735/X sky130_fd_sc_hd__xor2_1
XFILLER_61_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1746 U$$924/A1 U$$1746/A2 U$$789/A1 U$$1746/B2 VGND VGND VPWR VPWR U$$1747/A sky130_fd_sc_hd__a22o_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1757 U$$1757/A U$$1765/B VGND VGND VPWR VPWR U$$1757/X sky130_fd_sc_hd__xor2_1
XFILLER_199_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1768 U$$2316/A1 U$$1770/A2 U$$948/A1 U$$1770/B2 VGND VGND VPWR VPWR U$$1769/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1779 U$$1779/A U$$1779/B VGND VGND VPWR VPWR U$$1779/X sky130_fd_sc_hd__xor2_1
XFILLER_30_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_274 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_318_ _326_/CLK _318_/D VGND VGND VPWR VPWR _318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput12 a[1] VGND VGND VPWR VPWR U$$136/A sky130_fd_sc_hd__buf_6
Xinput23 a[2] VGND VGND VPWR VPWR U$$138/A sky130_fd_sc_hd__clkbuf_4
Xinput34 a[3] VGND VGND VPWR VPWR U$$274/A sky130_fd_sc_hd__buf_6
X_249_ _394_/CLK _249_/D VGND VGND VPWR VPWR _249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_554 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput45 a[4] VGND VGND VPWR VPWR U$$275/A sky130_fd_sc_hd__buf_2
XFILLER_122_1074 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput56 a[5] VGND VGND VPWR VPWR U$$410/A sky130_fd_sc_hd__buf_6
XFILLER_183_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput67 b[11] VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__buf_12
XFILLER_171_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput78 b[21] VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__buf_8
XFILLER_6_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput89 b[31] VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__buf_6
XFILLER_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_62_2 dadda_fa_2_62_2/A dadda_fa_2_62_2/B dadda_fa_2_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/A dadda_fa_3_62_3/A sky130_fd_sc_hd__fa_1
Xrepeater602 U$$1637/A2 VGND VGND VPWR VPWR U$$1635/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$409 final_adder.U$$408/B final_adder.U$$287/X final_adder.U$$283/X
+ VGND VGND VPWR VPWR final_adder.U$$409/X sky130_fd_sc_hd__a21o_1
Xrepeater613 U$$259/A2 VGND VGND VPWR VPWR U$$257/A2 sky130_fd_sc_hd__buf_6
XFILLER_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater624 U$$1361/A2 VGND VGND VPWR VPWR U$$1311/A2 sky130_fd_sc_hd__buf_4
XFILLER_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_55_1 dadda_fa_2_55_1/A dadda_fa_2_55_1/B dadda_fa_2_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_0/CIN dadda_fa_3_55_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater635 U$$1222/A2 VGND VGND VPWR VPWR U$$1190/A2 sky130_fd_sc_hd__buf_8
XFILLER_38_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater646 U$$1093/B2 VGND VGND VPWR VPWR U$$1083/B2 sky130_fd_sc_hd__buf_4
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater657 U$$690/X VGND VGND VPWR VPWR U$$793/B2 sky130_fd_sc_hd__buf_12
XU$$4350 U$$4350/A U$$4354/B VGND VGND VPWR VPWR U$$4350/X sky130_fd_sc_hd__xor2_1
Xrepeater668 U$$668/B2 VGND VGND VPWR VPWR U$$678/B2 sky130_fd_sc_hd__buf_6
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_32_0 dadda_fa_5_32_0/A dadda_fa_5_32_0/B dadda_fa_5_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_33_0/A dadda_fa_6_32_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater679 U$$537/B2 VGND VGND VPWR VPWR U$$491/B2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_48_0 U$$3162/X U$$3295/X U$$3321/B VGND VGND VPWR VPWR dadda_fa_3_49_0/B
+ dadda_fa_3_48_2/B sky130_fd_sc_hd__fa_1
XFILLER_168_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4361 U$$4498/A1 U$$4361/A2 U$$4361/B1 U$$4361/B2 VGND VGND VPWR VPWR U$$4362/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4372 U$$4372/A input60/X VGND VGND VPWR VPWR U$$4372/X sky130_fd_sc_hd__xor2_1
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4383 U$$4384/A VGND VGND VPWR VPWR U$$4383/Y sky130_fd_sc_hd__inv_1
XFILLER_80_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4394 U$$4394/A1 U$$4388/X U$$4396/A1 U$$4432/B2 VGND VGND VPWR VPWR U$$4395/A
+ sky130_fd_sc_hd__a22o_1
XU$$3660 U$$4343/B1 U$$3660/A2 U$$4210/A1 U$$3660/B2 VGND VGND VPWR VPWR U$$3661/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3671 U$$3671/A U$$3698/A VGND VGND VPWR VPWR U$$3671/X sky130_fd_sc_hd__xor2_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3682 U$$4365/B1 U$$3686/A2 U$$4095/A1 U$$3686/B2 VGND VGND VPWR VPWR U$$3683/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3693 U$$3693/A U$$3698/A VGND VGND VPWR VPWR U$$3693/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_17_clk clkbuf_3_1_0_clk/X VGND VGND VPWR VPWR _358_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$2970 U$$2970/A U$$2978/B VGND VGND VPWR VPWR U$$2970/X sky130_fd_sc_hd__xor2_1
XFILLER_209_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_9_1 input256/X dadda_fa_5_9_1/B dadda_ha_4_9_0/SUM VGND VGND VPWR VPWR
+ dadda_fa_6_10_0/B dadda_fa_7_9_0/A sky130_fd_sc_hd__fa_1
XFILLER_40_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2981 U$$3116/B1 U$$2985/A2 U$$2981/B1 U$$2985/B2 VGND VGND VPWR VPWR U$$2982/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2992 U$$2992/A U$$2996/B VGND VGND VPWR VPWR U$$2992/X sky130_fd_sc_hd__xor2_1
XFILLER_33_482 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_77_2 dadda_fa_4_77_2/A dadda_fa_4_77_2/B dadda_fa_4_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_78_0/CIN dadda_fa_5_77_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_161_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_47_0 dadda_fa_7_47_0/A dadda_fa_7_47_0/B dadda_fa_7_47_0/CIN VGND VGND
+ VPWR VPWR _344_/D _215_/D sky130_fd_sc_hd__fa_2
XFILLER_48_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$921 final_adder.U$$150/A final_adder.U$$859/X final_adder.U$$921/B1
+ VGND VGND VPWR VPWR final_adder.U$$921/X sky130_fd_sc_hd__a21o_1
XTAP_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$943 final_adder.U$$172/A final_adder.U$$881/X final_adder.U$$943/B1
+ VGND VGND VPWR VPWR final_adder.U$$943/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_0 U$$107/X U$$240/X U$$373/X VGND VGND VPWR VPWR dadda_fa_2_51_0/B
+ dadda_fa_2_50_3/B sky130_fd_sc_hd__fa_1
XFILLER_112_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$965 final_adder.U$$194/A final_adder.U$$807/X final_adder.U$$965/B1
+ VGND VGND VPWR VPWR final_adder.U$$965/X sky130_fd_sc_hd__a21o_1
XU$$804 U$$804/A U$$808/B VGND VGND VPWR VPWR U$$804/X sky130_fd_sc_hd__xor2_1
XFILLER_17_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$815 U$$950/B1 U$$689/X U$$954/A1 U$$690/X VGND VGND VPWR VPWR U$$816/A sky130_fd_sc_hd__a22o_1
XFILLER_95_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$987 final_adder.U$$216/A final_adder.U$$829/X final_adder.U$$987/B1
+ VGND VGND VPWR VPWR final_adder.U$$987/X sky130_fd_sc_hd__a21o_1
XU$$826 U$$824/Y input4/X input3/X U$$825/X U$$822/Y VGND VGND VPWR VPWR U$$826/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_71_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$837 U$$837/A U$$847/B VGND VGND VPWR VPWR U$$837/X sky130_fd_sc_hd__xor2_1
XFILLER_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$848 U$$983/B1 U$$872/A2 U$$850/A1 U$$872/B2 VGND VGND VPWR VPWR U$$849/A sky130_fd_sc_hd__a22o_1
XU$$859 U$$859/A U$$929/B VGND VGND VPWR VPWR U$$859/X sky130_fd_sc_hd__xor2_1
XFILLER_71_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1009 U$$598/A1 U$$997/A2 U$$598/B1 U$$997/B2 VGND VGND VPWR VPWR U$$1010/A sky130_fd_sc_hd__a22o_1
XFILLER_83_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_476 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_980 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1704 U$$3102/B1 VGND VGND VPWR VPWR U$$2282/A1 sky130_fd_sc_hd__buf_6
XFILLER_138_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4491_1822 VGND VGND VPWR VPWR U$$4491_1822/HI U$$4491/B sky130_fd_sc_hd__conb_1
XFILLER_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_72_1 dadda_fa_3_72_1/A dadda_fa_3_72_1/B dadda_fa_3_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_0/CIN dadda_fa_4_72_2/A sky130_fd_sc_hd__fa_1
XFILLER_140_549 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_65_0 dadda_fa_3_65_0/A dadda_fa_3_65_0/B dadda_fa_3_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_0/B dadda_fa_4_65_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_26_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2200 U$$2609/B1 U$$2252/A2 U$$2202/A1 U$$2252/B2 VGND VGND VPWR VPWR U$$2201/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2211 U$$2211/A U$$2227/B VGND VGND VPWR VPWR U$$2211/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_101_1 dadda_fa_4_101_1/A dadda_fa_4_101_1/B dadda_fa_4_101_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/B dadda_fa_5_101_1/B sky130_fd_sc_hd__fa_1
XU$$2222 U$$2357/B1 U$$2272/A2 U$$3594/A1 U$$2272/B2 VGND VGND VPWR VPWR U$$2223/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2233 U$$2233/A U$$2253/B VGND VGND VPWR VPWR U$$2233/X sky130_fd_sc_hd__xor2_1
XU$$2244 U$$3749/B1 U$$2284/A2 U$$3614/B1 U$$2284/B2 VGND VGND VPWR VPWR U$$2245/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1510 U$$1644/A U$$1510/B VGND VGND VPWR VPWR U$$1510/X sky130_fd_sc_hd__and2_1
XU$$2255 U$$2255/A U$$2303/B VGND VGND VPWR VPWR U$$2255/X sky130_fd_sc_hd__xor2_1
XU$$1521 U$$2343/A1 U$$1545/A2 U$$1932/B1 U$$1545/B2 VGND VGND VPWR VPWR U$$1522/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2266 U$$3499/A1 U$$2308/A2 U$$896/B1 U$$2308/B2 VGND VGND VPWR VPWR U$$2267/A
+ sky130_fd_sc_hd__a22o_1
XU$$2277 U$$2277/A U$$2303/B VGND VGND VPWR VPWR U$$2277/X sky130_fd_sc_hd__xor2_1
XFILLER_62_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1532 U$$1532/A U$$1546/B VGND VGND VPWR VPWR U$$1532/X sky130_fd_sc_hd__xor2_1
XU$$2288 U$$3245/B1 U$$2326/A2 U$$4480/B1 U$$2326/B2 VGND VGND VPWR VPWR U$$2289/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1543 U$$995/A1 U$$1545/A2 U$$997/A1 U$$1545/B2 VGND VGND VPWR VPWR U$$1544/A sky130_fd_sc_hd__a22o_1
XU$$1554 U$$1554/A U$$1558/B VGND VGND VPWR VPWR U$$1554/X sky130_fd_sc_hd__xor2_1
XU$$2299 U$$2299/A input27/X VGND VGND VPWR VPWR U$$2299/X sky130_fd_sc_hd__xor2_1
XU$$1565 U$$741/B1 U$$1591/A2 U$$745/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1566/A sky130_fd_sc_hd__a22o_1
XFILLER_203_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1576 U$$1576/A U$$1620/B VGND VGND VPWR VPWR U$$1576/X sky130_fd_sc_hd__xor2_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1587 U$$80/A1 U$$1621/A2 U$$2683/B1 U$$1621/B2 VGND VGND VPWR VPWR U$$1588/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_7_122_0 dadda_fa_7_122_0/A dadda_fa_7_122_0/B dadda_fa_7_122_0/CIN VGND
+ VGND VPWR VPWR _419_/D _290_/D sky130_fd_sc_hd__fa_1
XFILLER_176_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1598 U$$1598/A U$$1608/B VGND VGND VPWR VPWR U$$1598/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_496 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_87_1 dadda_fa_5_87_1/A dadda_fa_5_87_1/B dadda_fa_5_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_88_0/B dadda_fa_7_87_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_3_112_0_1866 VGND VGND VPWR VPWR dadda_fa_3_112_0/A dadda_fa_3_112_0_1866/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_171_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _323_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_103_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_79_8 U$$4288/X U$$4421/X input233/X VGND VGND VPWR VPWR dadda_fa_2_80_3/A
+ dadda_fa_3_79_0/A sky130_fd_sc_hd__fa_1
XFILLER_112_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$206 final_adder.U$$206/A final_adder.U$$206/B VGND VGND VPWR VPWR
+ final_adder.U$$334/B sky130_fd_sc_hd__and2_1
Xrepeater410 U$$652/A2 VGND VGND VPWR VPWR U$$578/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$217 final_adder.U$$216/B final_adder.U$$987/B1 final_adder.U$$217/B1
+ VGND VGND VPWR VPWR final_adder.U$$217/X sky130_fd_sc_hd__a21o_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater421 U$$4373/A2 VGND VGND VPWR VPWR U$$4369/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$228 final_adder.U$$228/A final_adder.U$$228/B VGND VGND VPWR VPWR
+ final_adder.U$$356/B sky130_fd_sc_hd__and2_1
Xrepeater432 U$$4176/A2 VGND VGND VPWR VPWR U$$4164/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$239 final_adder.U$$238/B final_adder.U$$239/A2 final_adder.U$$239/B1
+ VGND VGND VPWR VPWR final_adder.U$$239/X sky130_fd_sc_hd__a21o_1
Xrepeater443 U$$134/A2 VGND VGND VPWR VPWR U$$80/A2 sky130_fd_sc_hd__buf_6
XFILLER_100_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater454 U$$3977/X VGND VGND VPWR VPWR U$$4107/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater465 U$$3819/A2 VGND VGND VPWR VPWR U$$3813/A2 sky130_fd_sc_hd__buf_6
XFILLER_66_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater476 U$$3644/A2 VGND VGND VPWR VPWR U$$3696/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater487 U$$3292/X VGND VGND VPWR VPWR U$$3374/A2 sky130_fd_sc_hd__buf_6
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater498 U$$3155/X VGND VGND VPWR VPWR U$$3255/A2 sky130_fd_sc_hd__buf_4
XU$$4180 input89/X U$$4238/A2 input90/X U$$4238/B2 VGND VGND VPWR VPWR U$$4181/A sky130_fd_sc_hd__a22o_1
XFILLER_93_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4191 U$$4191/A U$$4211/B VGND VGND VPWR VPWR U$$4191/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3490 U$$3490/A U$$3490/B VGND VGND VPWR VPWR U$$3490/X sky130_fd_sc_hd__xor2_1
XFILLER_81_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_524 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_82_0 dadda_fa_4_82_0/A dadda_fa_4_82_0/B dadda_fa_4_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/A dadda_fa_5_82_1/A sky130_fd_sc_hd__fa_1
XFILLER_175_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_103_3 dadda_fa_3_103_3/A dadda_fa_3_103_3/B dadda_fa_3_103_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_104_1/B dadda_fa_4_103_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_175_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_579 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_868 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput202 c[50] VGND VGND VPWR VPWR input202/X sky130_fd_sc_hd__buf_2
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput213 c[60] VGND VGND VPWR VPWR input213/X sky130_fd_sc_hd__clkbuf_2
Xinput224 c[70] VGND VGND VPWR VPWR input224/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput235 c[80] VGND VGND VPWR VPWR input235/X sky130_fd_sc_hd__buf_2
XFILLER_88_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput246 c[90] VGND VGND VPWR VPWR input246/X sky130_fd_sc_hd__buf_2
XFILLER_75_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_338 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$740 final_adder.U$$772/B final_adder.U$$740/B VGND VGND VPWR VPWR
+ final_adder.U$$740/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$751 final_adder.U$$750/B final_adder.U$$671/X final_adder.U$$639/X
+ VGND VGND VPWR VPWR final_adder.U$$751/X sky130_fd_sc_hd__a21o_1
XFILLER_25_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$762 final_adder.U$$794/B final_adder.U$$762/B VGND VGND VPWR VPWR
+ final_adder.U$$762/X sky130_fd_sc_hd__and2_1
XTAP_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$601 U$$601/A U$$617/B VGND VGND VPWR VPWR U$$601/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$773 final_adder.U$$772/B final_adder.U$$693/X final_adder.U$$661/X
+ VGND VGND VPWR VPWR final_adder.U$$773/X sky130_fd_sc_hd__a21o_1
XTAP_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$612 U$$64/A1 U$$616/A2 U$$66/A1 U$$616/B2 VGND VGND VPWR VPWR U$$613/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$784 final_adder.U$$784/A final_adder.U$$784/B VGND VGND VPWR VPWR
+ final_adder.U$$784/X sky130_fd_sc_hd__and2_1
XFILLER_1_1028 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$623 U$$623/A U$$625/B VGND VGND VPWR VPWR U$$623/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$795 final_adder.U$$794/B final_adder.U$$715/X final_adder.U$$683/X
+ VGND VGND VPWR VPWR final_adder.U$$795/X sky130_fd_sc_hd__a21o_1
XFILLER_17_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$634 U$$84/B1 U$$636/A2 U$$910/A1 U$$636/B2 VGND VGND VPWR VPWR U$$635/A sky130_fd_sc_hd__a22o_1
XU$$645 U$$645/A U$$651/B VGND VGND VPWR VPWR U$$645/X sky130_fd_sc_hd__xor2_1
XFILLER_44_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$656 U$$930/A1 U$$678/A2 U$$930/B1 U$$678/B2 VGND VGND VPWR VPWR U$$657/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$667 U$$667/A U$$673/B VGND VGND VPWR VPWR U$$667/X sky130_fd_sc_hd__xor2_1
XFILLER_44_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$678 U$$950/B1 U$$678/A2 U$$678/B1 U$$678/B2 VGND VGND VPWR VPWR U$$679/A sky130_fd_sc_hd__a22o_1
XU$$689 U$$687/Y input2/X U$$685/A U$$688/X U$$685/Y VGND VGND VPWR VPWR U$$689/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_32_728 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_97_0 dadda_fa_6_97_0/A dadda_fa_6_97_0/B dadda_fa_6_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_98_0/B dadda_fa_7_97_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_200_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_438 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1501 U$$4379/A1 VGND VGND VPWR VPWR U$$4516/A1 sky130_fd_sc_hd__buf_6
Xrepeater1512 input122/X VGND VGND VPWR VPWR U$$4240/A1 sky130_fd_sc_hd__buf_6
Xrepeater1523 U$$3032/A1 VGND VGND VPWR VPWR U$$18/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1534 U$$127/B VGND VGND VPWR VPWR U$$111/B sky130_fd_sc_hd__buf_8
Xrepeater1545 input119/X VGND VGND VPWR VPWR U$$3551/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1556 input117/X VGND VGND VPWR VPWR U$$3684/A1 sky130_fd_sc_hd__buf_4
XFILLER_181_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1567 U$$2449/A1 VGND VGND VPWR VPWR U$$2312/A1 sky130_fd_sc_hd__buf_8
XFILLER_119_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1578 input115/X VGND VGND VPWR VPWR U$$3817/A1 sky130_fd_sc_hd__buf_4
XFILLER_158_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1589 U$$2032/A1 VGND VGND VPWR VPWR U$$936/A1 sky130_fd_sc_hd__buf_4
XFILLER_165_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_33_5 U$$2068/X U$$2201/X VGND VGND VPWR VPWR dadda_fa_3_34_2/A dadda_fa_4_33_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_79_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_32_3 U$$1268/X U$$1401/X U$$1534/X VGND VGND VPWR VPWR dadda_fa_3_33_1/B
+ dadda_fa_3_32_3/B sky130_fd_sc_hd__fa_1
XU$$2030 U$$2715/A1 U$$2046/A2 U$$2032/A1 U$$2046/B2 VGND VGND VPWR VPWR U$$2031/A
+ sky130_fd_sc_hd__a22o_1
XU$$2041 U$$2041/A U$$2043/B VGND VGND VPWR VPWR U$$2041/X sky130_fd_sc_hd__xor2_1
XU$$2052 U$$3283/B1 U$$2052/A2 U$$2052/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2053/A
+ sky130_fd_sc_hd__a22o_1
XU$$2063 U$$2198/B1 U$$2093/A2 U$$2063/B1 U$$2093/B2 VGND VGND VPWR VPWR U$$2064/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2074 U$$2074/A U$$2100/B VGND VGND VPWR VPWR U$$2074/X sky130_fd_sc_hd__xor2_1
XU$$1340 U$$1340/A U$$1370/A VGND VGND VPWR VPWR U$$1340/X sky130_fd_sc_hd__xor2_1
XFILLER_90_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2085 U$$2357/B1 U$$2091/A2 U$$3594/A1 U$$2091/B2 VGND VGND VPWR VPWR U$$2086/A
+ sky130_fd_sc_hd__a22o_1
XU$$2096 U$$2096/A U$$2100/B VGND VGND VPWR VPWR U$$2096/X sky130_fd_sc_hd__xor2_1
XU$$1351 U$$527/B1 U$$1361/A2 U$$2449/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1352/A
+ sky130_fd_sc_hd__a22o_1
XU$$1362 U$$1362/A U$$1366/B VGND VGND VPWR VPWR U$$1362/X sky130_fd_sc_hd__xor2_1
XFILLER_204_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1373 U$$1507/A U$$1373/B VGND VGND VPWR VPWR U$$1373/X sky130_fd_sc_hd__and2_1
XFILLER_50_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1384 U$$2069/A1 U$$1404/A2 U$$1932/B1 U$$1404/B2 VGND VGND VPWR VPWR U$$1385/A
+ sky130_fd_sc_hd__a22o_1
XU$$1395 U$$1395/A U$$1399/B VGND VGND VPWR VPWR U$$1395/X sky130_fd_sc_hd__xor2_1
XFILLER_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_77_5 U$$3353/X U$$3486/X U$$3619/X VGND VGND VPWR VPWR dadda_fa_2_78_2/A
+ dadda_fa_2_77_5/A sky130_fd_sc_hd__fa_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$80 _376_/Q _248_/Q VGND VGND VPWR VPWR final_adder.U$$945/B1 final_adder.U$$174/A
+ sky130_fd_sc_hd__ha_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$91 _387_/Q _259_/Q VGND VGND VPWR VPWR final_adder.U$$165/B1 final_adder.U$$164/B
+ sky130_fd_sc_hd__ha_1
XFILLER_186_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_101_0 U$$4199/X U$$4332/X U$$4465/X VGND VGND VPWR VPWR dadda_fa_4_102_0/B
+ dadda_fa_4_101_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_108_899 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_65_3 U$$1334/X U$$1467/X U$$1600/X VGND VGND VPWR VPWR dadda_fa_1_66_6/B
+ dadda_fa_1_65_8/B sky130_fd_sc_hd__fa_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_42_2 dadda_fa_3_42_2/A dadda_fa_3_42_2/B dadda_fa_3_42_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_1/A dadda_fa_4_42_2/B sky130_fd_sc_hd__fa_1
XFILLER_97_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_58_2 U$$921/X U$$1054/X U$$1187/X VGND VGND VPWR VPWR dadda_fa_1_59_7/B
+ dadda_fa_1_58_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$570 final_adder.U$$578/B final_adder.U$$570/B VGND VGND VPWR VPWR
+ final_adder.U$$690/B sky130_fd_sc_hd__and2_1
XTAP_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_35_1 dadda_fa_3_35_1/A dadda_fa_3_35_1/B dadda_fa_3_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_0/CIN dadda_fa_4_35_2/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$581 final_adder.U$$580/B final_adder.U$$465/X final_adder.U$$457/X
+ VGND VGND VPWR VPWR final_adder.U$$581/X sky130_fd_sc_hd__a21o_1
XTAP_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$420 U$$420/A U$$436/B VGND VGND VPWR VPWR U$$420/X sky130_fd_sc_hd__xor2_1
XTAP_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$592 final_adder.U$$600/B final_adder.U$$592/B VGND VGND VPWR VPWR
+ final_adder.U$$712/B sky130_fd_sc_hd__and2_1
XU$$431 U$$431/A1 U$$515/A2 U$$842/B1 U$$515/B2 VGND VGND VPWR VPWR U$$432/A sky130_fd_sc_hd__a22o_1
XTAP_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$442 U$$442/A U$$474/B VGND VGND VPWR VPWR U$$442/X sky130_fd_sc_hd__xor2_1
XFILLER_44_330 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_12_0 dadda_fa_6_12_0/A dadda_fa_6_12_0/B dadda_fa_6_12_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_13_0/B dadda_fa_7_12_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$453 U$$42/A1 U$$473/A2 U$$866/A1 U$$473/B2 VGND VGND VPWR VPWR U$$454/A sky130_fd_sc_hd__a22o_1
XTAP_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_28_0 U$$1526/X U$$1659/X U$$1792/X VGND VGND VPWR VPWR dadda_fa_4_29_0/B
+ dadda_fa_4_28_1/CIN sky130_fd_sc_hd__fa_1
XU$$464 U$$464/A U$$484/B VGND VGND VPWR VPWR U$$464/X sky130_fd_sc_hd__xor2_1
XFILLER_204_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$475 U$$610/B1 U$$527/A2 U$$477/A1 U$$527/B2 VGND VGND VPWR VPWR U$$476/A sky130_fd_sc_hd__a22o_1
XU$$486 U$$486/A U$$492/B VGND VGND VPWR VPWR U$$486/X sky130_fd_sc_hd__xor2_1
XFILLER_44_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$497 U$$86/A1 U$$537/A2 U$$88/A1 U$$537/B2 VGND VGND VPWR VPWR U$$498/A sky130_fd_sc_hd__a22o_1
XFILLER_204_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1320 U$$3288/A VGND VGND VPWR VPWR U$$3244/B sky130_fd_sc_hd__buf_8
Xdadda_fa_2_94_5 dadda_fa_2_94_5/A dadda_fa_2_94_5/B dadda_fa_2_94_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_95_2/A dadda_fa_4_94_0/A sky130_fd_sc_hd__fa_1
Xrepeater1331 U$$2950/B VGND VGND VPWR VPWR U$$2922/B sky130_fd_sc_hd__buf_8
XFILLER_172_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1342 U$$2825/B VGND VGND VPWR VPWR U$$2817/B sky130_fd_sc_hd__buf_8
XFILLER_99_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1353 U$$244/B VGND VGND VPWR VPWR U$$212/B sky130_fd_sc_hd__buf_6
XFILLER_181_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_87_4 dadda_fa_2_87_4/A dadda_fa_2_87_4/B dadda_fa_2_87_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_1/CIN dadda_fa_3_87_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1364 input33/X VGND VGND VPWR VPWR U$$2710/B sky130_fd_sc_hd__buf_8
XFILLER_114_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1375 U$$784/B VGND VGND VPWR VPWR U$$712/B sky130_fd_sc_hd__buf_6
XFILLER_113_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1386 U$$2446/B VGND VGND VPWR VPWR U$$2426/B sky130_fd_sc_hd__buf_8
XFILLER_99_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1397 U$$2317/B VGND VGND VPWR VPWR U$$2328/A sky130_fd_sc_hd__buf_6
XFILLER_114_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_24_1 U$$454/X U$$587/X VGND VGND VPWR VPWR dadda_fa_3_25_3/B dadda_fa_4_24_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_55_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_30_0 U$$67/X U$$200/X U$$333/X VGND VGND VPWR VPWR dadda_fa_3_31_1/A dadda_fa_3_30_2/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_39_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_103_2 U$$3538/X U$$3671/X U$$3804/X VGND VGND VPWR VPWR dadda_fa_3_104_3/A
+ dadda_fa_4_103_0/A sky130_fd_sc_hd__fa_1
XFILLER_165_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1170 U$$74/A1 U$$1174/A2 U$$1446/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1171/A sky130_fd_sc_hd__a22o_1
XU$$1181 U$$1181/A U$$1223/B VGND VGND VPWR VPWR U$$1181/X sky130_fd_sc_hd__xor2_1
XU$$1192 U$$96/A1 U$$1204/A2 U$$98/A1 U$$1204/B2 VGND VGND VPWR VPWR U$$1193/A sky130_fd_sc_hd__a22o_1
XFILLER_148_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_117_0 dadda_fa_5_117_0/A dadda_fa_5_117_0/B dadda_fa_5_117_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_118_0/A dadda_fa_6_117_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_15_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_983 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_82_3 U$$2432/X U$$2565/X U$$2698/X VGND VGND VPWR VPWR dadda_fa_2_83_2/B
+ dadda_fa_2_82_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1059 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_75_2 U$$2418/X U$$2551/X U$$2684/X VGND VGND VPWR VPWR dadda_fa_2_76_1/A
+ dadda_fa_2_75_4/A sky130_fd_sc_hd__fa_1
XFILLER_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_52_1 dadda_fa_4_52_1/A dadda_fa_4_52_1/B dadda_fa_4_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/B dadda_fa_5_52_1/B sky130_fd_sc_hd__fa_1
XFILLER_59_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_68_1 U$$2936/X U$$3069/X U$$3202/X VGND VGND VPWR VPWR dadda_fa_2_69_0/CIN
+ dadda_fa_2_68_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_45_0 dadda_fa_4_45_0/A dadda_fa_4_45_0/B dadda_fa_4_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/A dadda_fa_5_45_1/A sky130_fd_sc_hd__fa_1
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _384_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_115 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _390_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_420_ _420_/CLK _420_/D VGND VGND VPWR VPWR _420_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_137 input168/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 input65/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_159 U$$2691/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_351_ _351_/CLK _351_/D VGND VGND VPWR VPWR _351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_1117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_282_ _420_/CLK _282_/D VGND VGND VPWR VPWR _282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_97_3 dadda_fa_3_97_3/A dadda_fa_3_97_3/B dadda_fa_3_97_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_98_1/B dadda_fa_4_97_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_30_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_0_70_1 U$$812/X U$$945/X U$$1078/X VGND VGND VPWR VPWR dadda_fa_1_71_6/CIN
+ dadda_fa_1_70_8/A sky130_fd_sc_hd__fa_1
XFILLER_122_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_0_63_0 U$$133/X U$$266/X U$$399/X VGND VGND VPWR VPWR dadda_fa_1_64_5/B
+ dadda_fa_1_63_7/B sky130_fd_sc_hd__fa_1
XTAP_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_943 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$250 U$$250/A U$$260/B VGND VGND VPWR VPWR U$$250/X sky130_fd_sc_hd__xor2_1
XTAP_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$261 U$$944/B1 U$$141/X U$$674/A1 U$$142/X VGND VGND VPWR VPWR U$$262/A sky130_fd_sc_hd__a22o_1
XU$$272 U$$272/A U$$272/B VGND VGND VPWR VPWR U$$272/X sky130_fd_sc_hd__xor2_2
XU$$283 U$$283/A U$$317/B VGND VGND VPWR VPWR U$$283/X sky130_fd_sc_hd__xor2_1
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$294 U$$20/A1 U$$302/A2 U$$22/A1 U$$302/B2 VGND VGND VPWR VPWR U$$295/A sky130_fd_sc_hd__a22o_1
XFILLER_44_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$0 U$$0/A VGND VGND VPWR VPWR U$$0/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$8 _304_/Q _176_/Q VGND VGND VPWR VPWR final_adder.U$$8/COUT final_adder.U$$8/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_173_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput303 output303/A VGND VGND VPWR VPWR o[26] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_2 U$$3782/X U$$3915/X U$$4048/X VGND VGND VPWR VPWR dadda_fa_3_93_1/A
+ dadda_fa_3_92_3/A sky130_fd_sc_hd__fa_1
Xoutput314 output314/A VGND VGND VPWR VPWR o[36] sky130_fd_sc_hd__buf_2
XFILLER_195_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput325 output325/A VGND VGND VPWR VPWR o[46] sky130_fd_sc_hd__buf_2
Xoutput336 output336/A VGND VGND VPWR VPWR o[56] sky130_fd_sc_hd__buf_2
Xrepeater1150 U$$4144/B1 VGND VGND VPWR VPWR U$$4009/A1 sky130_fd_sc_hd__buf_8
Xoutput347 output347/A VGND VGND VPWR VPWR o[66] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_85_1 U$$4300/X U$$4433/X input240/X VGND VGND VPWR VPWR dadda_fa_3_86_0/CIN
+ dadda_fa_3_85_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater1161 U$$962/A VGND VGND VPWR VPWR U$$1076/B sky130_fd_sc_hd__buf_6
Xoutput358 output358/A VGND VGND VPWR VPWR o[76] sky130_fd_sc_hd__buf_2
Xrepeater1172 U$$3183/A1 VGND VGND VPWR VPWR U$$854/A1 sky130_fd_sc_hd__buf_4
Xoutput369 output369/A VGND VGND VPWR VPWR o[86] sky130_fd_sc_hd__buf_2
Xrepeater1183 input67/X VGND VGND VPWR VPWR U$$578/A1 sky130_fd_sc_hd__buf_4
Xrepeater1194 U$$4275/A1 VGND VGND VPWR VPWR U$$4273/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_62_0 dadda_fa_5_62_0/A dadda_fa_5_62_0/B dadda_fa_5_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_63_0/A dadda_fa_6_62_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_78_0 dadda_fa_2_78_0/A dadda_fa_2_78_0/B dadda_fa_2_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_0/B dadda_fa_3_78_2/B sky130_fd_sc_hd__fa_1
XFILLER_142_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_61_8 dadda_fa_1_61_8/A dadda_fa_1_61_8/B dadda_fa_1_61_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_62_3/A dadda_fa_3_61_0/A sky130_fd_sc_hd__fa_2
XFILLER_206_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_54_7 U$$3573/X U$$3706/X U$$3794/B VGND VGND VPWR VPWR dadda_fa_2_55_2/CIN
+ dadda_fa_2_54_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_1112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_831 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_77_0 dadda_fa_7_77_0/A dadda_fa_7_77_0/B dadda_fa_7_77_0/CIN VGND VGND
+ VPWR VPWR _374_/D _245_/D sky130_fd_sc_hd__fa_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_80_0 dadda_fa_1_80_0/A U$$1231/X U$$1364/X VGND VGND VPWR VPWR dadda_fa_2_81_0/CIN
+ dadda_fa_2_80_3/B sky130_fd_sc_hd__fa_1
XFILLER_78_506 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4009 U$$4009/A1 U$$4043/A2 U$$4422/A1 U$$4043/B2 VGND VGND VPWR VPWR U$$4010/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_926 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3308 U$$431/A1 U$$3394/A2 input126/X U$$3394/B2 VGND VGND VPWR VPWR U$$3309/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3319 U$$3319/A U$$3321/B VGND VGND VPWR VPWR U$$3319/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2607 U$$2605/Y input32/X input31/X U$$2606/X U$$2603/Y VGND VGND VPWR VPWR U$$2607/X
+ sky130_fd_sc_hd__a32o_4
XU$$2618 U$$2618/A U$$2624/B VGND VGND VPWR VPWR U$$2618/X sky130_fd_sc_hd__xor2_1
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2629 U$$3451/A1 U$$2653/A2 U$$711/B1 U$$2653/B2 VGND VGND VPWR VPWR U$$2630/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1906 U$$1906/A U$$1912/B VGND VGND VPWR VPWR U$$1906/X sky130_fd_sc_hd__xor2_1
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1917 U$$1917/A VGND VGND VPWR VPWR U$$1917/Y sky130_fd_sc_hd__inv_1
XFILLER_148_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1928 U$$2063/B1 U$$1990/A2 U$$2065/B1 U$$1990/B2 VGND VGND VPWR VPWR U$$1929/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_403_ _407_/CLK _403_/D VGND VGND VPWR VPWR _403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1939 U$$1939/A U$$1971/B VGND VGND VPWR VPWR U$$1939/X sky130_fd_sc_hd__xor2_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ _342_/CLK _334_/D VGND VGND VPWR VPWR _334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_265_ _394_/CLK _265_/D VGND VGND VPWR VPWR _265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_196_ _329_/CLK _196_/D VGND VGND VPWR VPWR _196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4455_1804 VGND VGND VPWR VPWR U$$4455_1804/HI U$$4455/B sky130_fd_sc_hd__conb_1
XFILLER_109_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_95_0 dadda_fa_3_95_0/A dadda_fa_3_95_0/B dadda_fa_3_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_0/B dadda_fa_4_95_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_183_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1098 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater806 U$$2197/X VGND VGND VPWR VPWR U$$2308/B2 sky130_fd_sc_hd__buf_4
XFILLER_42_1224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater817 U$$2149/B2 VGND VGND VPWR VPWR U$$2099/B2 sky130_fd_sc_hd__buf_4
Xrepeater828 U$$2040/B2 VGND VGND VPWR VPWR U$$1960/B2 sky130_fd_sc_hd__buf_4
Xrepeater839 U$$1736/B2 VGND VGND VPWR VPWR U$$1688/B2 sky130_fd_sc_hd__buf_4
XU$$4510 U$$4510/A1 U$$4388/X U$$4512/A1 U$$4512/B2 VGND VGND VPWR VPWR U$$4511/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_57_5 dadda_fa_2_57_5/A dadda_fa_2_57_5/B dadda_fa_2_57_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_58_2/A dadda_fa_4_57_0/A sky130_fd_sc_hd__fa_2
XFILLER_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$13 U$$13/A U$$9/B VGND VGND VPWR VPWR U$$13/X sky130_fd_sc_hd__xor2_1
XU$$24 U$$24/A1 U$$8/A2 U$$26/A1 U$$8/B2 VGND VGND VPWR VPWR U$$25/A sky130_fd_sc_hd__a22o_1
XU$$3820 U$$3820/A U$$3826/B VGND VGND VPWR VPWR U$$3820/X sky130_fd_sc_hd__xor2_1
XU$$35 U$$35/A U$$51/B VGND VGND VPWR VPWR U$$35/X sky130_fd_sc_hd__xor2_1
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3831 U$$4379/A1 U$$3833/A2 input124/X U$$3833/B2 VGND VGND VPWR VPWR U$$3832/A
+ sky130_fd_sc_hd__a22o_1
XU$$46 U$$46/A1 U$$50/A2 U$$48/A1 U$$50/B2 VGND VGND VPWR VPWR U$$47/A sky130_fd_sc_hd__a22o_1
XTAP_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3842 U$$3842/A1 U$$3926/A2 U$$3979/B1 U$$3926/B2 VGND VGND VPWR VPWR U$$3843/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$57 U$$57/A U$$85/B VGND VGND VPWR VPWR U$$57/X sky130_fd_sc_hd__xor2_1
XTAP_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3853 U$$3853/A U$$3875/B VGND VGND VPWR VPWR U$$3853/X sky130_fd_sc_hd__xor2_1
XU$$3864 U$$4273/B1 U$$3902/A2 U$$4275/B1 U$$3902/B2 VGND VGND VPWR VPWR U$$3865/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$68 U$$68/A1 U$$80/A2 U$$70/A1 U$$80/B2 VGND VGND VPWR VPWR U$$69/A sky130_fd_sc_hd__a22o_1
XU$$79 U$$79/A U$$81/B VGND VGND VPWR VPWR U$$79/X sky130_fd_sc_hd__xor2_1
XU$$3875 U$$3875/A U$$3875/B VGND VGND VPWR VPWR U$$3875/X sky130_fd_sc_hd__xor2_1
XU$$3886 U$$50/A1 U$$3970/A2 input79/X U$$3970/B2 VGND VGND VPWR VPWR U$$3887/A sky130_fd_sc_hd__a22o_1
XFILLER_206_773 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3897 U$$3897/A U$$3903/B VGND VGND VPWR VPWR U$$3897/X sky130_fd_sc_hd__xor2_1
XFILLER_205_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_15 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_26 _337_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_37 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_308 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_48 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_59 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_52_4 U$$1973/X U$$2106/X U$$2239/X VGND VGND VPWR VPWR dadda_fa_2_53_1/CIN
+ dadda_fa_2_52_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_49 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_45_3 U$$1294/X U$$1427/X U$$1560/X VGND VGND VPWR VPWR dadda_fa_2_46_3/A
+ dadda_fa_2_45_5/B sky130_fd_sc_hd__fa_1
XFILLER_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_22_2 dadda_fa_4_22_2/A dadda_fa_4_22_2/B dadda_fa_4_22_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_23_0/CIN dadda_fa_5_22_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_15_1 U$$702/X U$$835/X U$$968/X VGND VGND VPWR VPWR dadda_fa_5_16_0/B
+ dadda_fa_5_15_1/B sky130_fd_sc_hd__fa_1
XFILLER_145_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_675 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1007 final_adder.U$$236/A final_adder.U$$737/X final_adder.U$$237/A2
+ VGND VGND VPWR VPWR final_adder.U$$1043/B sky130_fd_sc_hd__a21o_1
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1029 final_adder.U$$5/SUM final_adder.U$$1029/B VGND VGND VPWR VPWR
+ output340/A sky130_fd_sc_hd__xor2_1
XFILLER_183_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4485_1819 VGND VGND VPWR VPWR U$$4485_1819/HI U$$4485/B sky130_fd_sc_hd__conb_1
XFILLER_87_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3105 U$$3105/A U$$3109/B VGND VGND VPWR VPWR U$$3105/X sky130_fd_sc_hd__xor2_1
XFILLER_47_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3116 U$$3116/A1 U$$3118/A2 U$$3116/B1 U$$3118/B2 VGND VGND VPWR VPWR U$$3117/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3127 U$$3127/A U$$3133/B VGND VGND VPWR VPWR U$$3127/X sky130_fd_sc_hd__xor2_1
XFILLER_207_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3138 U$$3684/B1 U$$3148/A2 U$$3551/A1 U$$3148/B2 VGND VGND VPWR VPWR U$$3139/A
+ sky130_fd_sc_hd__a22o_1
XU$$2404 U$$2404/A U$$2442/B VGND VGND VPWR VPWR U$$2404/X sky130_fd_sc_hd__xor2_1
XFILLER_74_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3149 U$$3149/A U$$3150/A VGND VGND VPWR VPWR U$$3149/X sky130_fd_sc_hd__xor2_1
XFILLER_35_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2415 U$$2415/A1 U$$2435/A2 U$$2415/B1 U$$2435/B2 VGND VGND VPWR VPWR U$$2416/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2426 U$$2426/A U$$2426/B VGND VGND VPWR VPWR U$$2426/X sky130_fd_sc_hd__xor2_1
XU$$2437 U$$2709/B1 U$$2333/X U$$2711/B1 U$$2334/X VGND VGND VPWR VPWR U$$2438/A sky130_fd_sc_hd__a22o_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2448 U$$2448/A U$$2454/B VGND VGND VPWR VPWR U$$2448/X sky130_fd_sc_hd__xor2_1
XFILLER_61_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1703 U$$1703/A U$$1707/B VGND VGND VPWR VPWR U$$1703/X sky130_fd_sc_hd__xor2_1
XU$$2459 U$$3281/A1 U$$2459/A2 U$$3281/B1 U$$2459/B2 VGND VGND VPWR VPWR U$$2460/A
+ sky130_fd_sc_hd__a22o_1
XU$$1714 U$$1714/A1 U$$1750/A2 U$$2949/A1 U$$1750/B2 VGND VGND VPWR VPWR U$$1715/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1725 U$$1725/A U$$1739/B VGND VGND VPWR VPWR U$$1725/X sky130_fd_sc_hd__xor2_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1736 U$$2967/B1 U$$1736/A2 U$$3108/A1 U$$1736/B2 VGND VGND VPWR VPWR U$$1737/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1747 U$$1747/A U$$1780/A VGND VGND VPWR VPWR U$$1747/X sky130_fd_sc_hd__xor2_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1758 U$$2717/A1 U$$1764/A2 U$$2582/A1 U$$1764/B2 VGND VGND VPWR VPWR U$$1759/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1769 U$$1769/A U$$1780/A VGND VGND VPWR VPWR U$$1769/X sky130_fd_sc_hd__xor2_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_317_ _327_/CLK _317_/D VGND VGND VPWR VPWR _317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 a[20] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput24 a[30] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
X_248_ _379_/CLK _248_/D VGND VGND VPWR VPWR _248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput35 a[40] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 a[50] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_566 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput57 a[60] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput68 b[12] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__buf_6
XFILLER_122_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_179_ _327_/CLK _179_/D VGND VGND VPWR VPWR _179_/Q sky130_fd_sc_hd__dfxtp_1
Xinput79 b[22] VGND VGND VPWR VPWR input79/X sky130_fd_sc_hd__buf_8
XFILLER_157_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_62_3 dadda_fa_2_62_3/A dadda_fa_2_62_3/B dadda_fa_2_62_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/B dadda_fa_3_62_3/B sky130_fd_sc_hd__fa_1
XFILLER_69_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater603 U$$1557/A2 VGND VGND VPWR VPWR U$$1545/A2 sky130_fd_sc_hd__buf_4
XFILLER_69_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater614 U$$141/X VGND VGND VPWR VPWR U$$259/A2 sky130_fd_sc_hd__buf_4
XFILLER_78_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater625 U$$1367/A2 VGND VGND VPWR VPWR U$$1361/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_55_2 dadda_fa_2_55_2/A dadda_fa_2_55_2/B dadda_fa_2_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/A dadda_fa_3_55_3/A sky130_fd_sc_hd__fa_1
Xrepeater636 U$$1100/X VGND VGND VPWR VPWR U$$1222/A2 sky130_fd_sc_hd__buf_6
Xrepeater647 U$$964/X VGND VGND VPWR VPWR U$$1093/B2 sky130_fd_sc_hd__buf_8
Xrepeater658 U$$749/B2 VGND VGND VPWR VPWR U$$739/B2 sky130_fd_sc_hd__buf_4
XU$$4340 U$$4340/A U$$4354/B VGND VGND VPWR VPWR U$$4340/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_32_1 dadda_fa_5_32_1/A dadda_fa_5_32_1/B dadda_fa_5_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_33_0/B dadda_fa_7_32_0/A sky130_fd_sc_hd__fa_1
XU$$4351 input107/X U$$4373/A2 input108/X U$$4373/B2 VGND VGND VPWR VPWR U$$4352/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater669 U$$553/X VGND VGND VPWR VPWR U$$668/B2 sky130_fd_sc_hd__buf_4
XU$$4362 U$$4362/A U$$4366/B VGND VGND VPWR VPWR U$$4362/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_48_1 input199/X dadda_fa_2_48_1/B dadda_fa_2_48_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_49_0/CIN dadda_fa_3_48_2/CIN sky130_fd_sc_hd__fa_1
XU$$4373 U$$4510/A1 U$$4373/A2 U$$4512/A1 U$$4373/B2 VGND VGND VPWR VPWR U$$4374/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4384 U$$4384/A VGND VGND VPWR VPWR U$$4384/Y sky130_fd_sc_hd__inv_1
XFILLER_38_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_25_0 dadda_fa_5_25_0/A dadda_fa_5_25_0/B dadda_fa_5_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_26_0/A dadda_fa_6_25_0/CIN sky130_fd_sc_hd__fa_1
XU$$3650 U$$4333/B1 U$$3686/A2 U$$3787/B1 U$$3686/B2 VGND VGND VPWR VPWR U$$3651/A
+ sky130_fd_sc_hd__a22o_1
XU$$4395 U$$4395/A U$$4395/B VGND VGND VPWR VPWR U$$4395/X sky130_fd_sc_hd__xor2_1
XU$$3661 U$$3661/A U$$3665/B VGND VGND VPWR VPWR U$$3661/X sky130_fd_sc_hd__xor2_1
XU$$3672 U$$3944/B1 U$$3680/A2 U$$3946/B1 U$$3680/B2 VGND VGND VPWR VPWR U$$3673/A
+ sky130_fd_sc_hd__a22o_1
XU$$3683 U$$3683/A U$$3683/B VGND VGND VPWR VPWR U$$3683/X sky130_fd_sc_hd__xor2_1
XFILLER_37_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3694 U$$4379/A1 U$$3696/A2 input124/X U$$3696/B2 VGND VGND VPWR VPWR U$$3695/A
+ sky130_fd_sc_hd__a22o_1
XU$$2960 U$$2960/A U$$3008/B VGND VGND VPWR VPWR U$$2960/X sky130_fd_sc_hd__xor2_1
XU$$2971 U$$3108/A1 U$$2977/A2 U$$3108/B1 U$$2979/B2 VGND VGND VPWR VPWR U$$2972/A
+ sky130_fd_sc_hd__a22o_1
XU$$2982 U$$2982/A U$$3008/B VGND VGND VPWR VPWR U$$2982/X sky130_fd_sc_hd__xor2_1
XU$$2993 U$$388/B1 U$$2995/A2 U$$3680/A1 U$$2995/B2 VGND VGND VPWR VPWR U$$2994/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_26 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_1_37_1 U$$480/X U$$613/X VGND VGND VPWR VPWR dadda_fa_2_38_5/A dadda_fa_3_37_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$911 final_adder.U$$140/A final_adder.U$$849/X final_adder.U$$911/B1
+ VGND VGND VPWR VPWR final_adder.U$$911/X sky130_fd_sc_hd__a21o_1
XTAP_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$933 final_adder.U$$162/A final_adder.U$$871/X final_adder.U$$933/B1
+ VGND VGND VPWR VPWR final_adder.U$$933/X sky130_fd_sc_hd__a21o_1
XTAP_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_50_1 U$$506/X U$$639/X U$$772/X VGND VGND VPWR VPWR dadda_fa_2_51_0/CIN
+ dadda_fa_2_50_3/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$955 final_adder.U$$184/A final_adder.U$$893/X final_adder.U$$955/B1
+ VGND VGND VPWR VPWR final_adder.U$$955/X sky130_fd_sc_hd__a21o_1
XFILLER_60_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$805 U$$940/B1 U$$805/A2 U$$807/A1 U$$805/B2 VGND VGND VPWR VPWR U$$806/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$977 final_adder.U$$206/A final_adder.U$$819/X final_adder.U$$977/B1
+ VGND VGND VPWR VPWR final_adder.U$$977/X sky130_fd_sc_hd__a21o_1
XFILLER_21_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$816 U$$816/A U$$821/A VGND VGND VPWR VPWR U$$816/X sky130_fd_sc_hd__xor2_1
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$827 U$$825/B input3/X input4/X U$$822/Y VGND VGND VPWR VPWR U$$827/X sky130_fd_sc_hd__a22o_4
Xdadda_fa_1_43_0 U$$93/X U$$226/X U$$359/X VGND VGND VPWR VPWR dadda_fa_2_44_2/CIN
+ dadda_fa_2_43_4/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$999 final_adder.U$$228/A final_adder.U$$729/X final_adder.U$$999/B1
+ VGND VGND VPWR VPWR final_adder.U$$999/X sky130_fd_sc_hd__a21o_1
XU$$838 U$$16/A1 U$$872/A2 U$$18/A1 U$$872/B2 VGND VGND VPWR VPWR U$$839/A sky130_fd_sc_hd__a22o_1
XFILLER_83_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$849 U$$849/A U$$877/B VGND VGND VPWR VPWR U$$849/X sky130_fd_sc_hd__xor2_1
XFILLER_56_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_915 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1705 U$$4335/B1 VGND VGND VPWR VPWR U$$3102/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_193_992 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_72_2 dadda_fa_3_72_2/A dadda_fa_3_72_2/B dadda_fa_3_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_1/A dadda_fa_4_72_2/B sky130_fd_sc_hd__fa_1
XFILLER_3_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_65_1 dadda_fa_3_65_1/A dadda_fa_3_65_1/B dadda_fa_3_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_0/CIN dadda_fa_4_65_2/A sky130_fd_sc_hd__fa_1
XFILLER_191_1095 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_42_0 dadda_fa_6_42_0/A dadda_fa_6_42_0/B dadda_fa_6_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_43_0/B dadda_fa_7_42_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_117_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_58_0 dadda_fa_3_58_0/A dadda_fa_3_58_0/B dadda_fa_3_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_0/B dadda_fa_4_58_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_208_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2201 U$$2201/A U$$2253/B VGND VGND VPWR VPWR U$$2201/X sky130_fd_sc_hd__xor2_1
XU$$2212 U$$2623/A1 U$$2226/A2 U$$2625/A1 U$$2226/B2 VGND VGND VPWR VPWR U$$2213/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_101_2 dadda_fa_4_101_2/A dadda_fa_4_101_2/B dadda_fa_4_101_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_102_0/CIN dadda_fa_5_101_1/CIN sky130_fd_sc_hd__fa_1
XU$$2223 U$$2223/A U$$2273/B VGND VGND VPWR VPWR U$$2223/X sky130_fd_sc_hd__xor2_1
XFILLER_62_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2234 U$$179/A1 U$$2284/A2 U$$44/A1 U$$2284/B2 VGND VGND VPWR VPWR U$$2235/A sky130_fd_sc_hd__a22o_1
XU$$2245 U$$2245/A U$$2285/B VGND VGND VPWR VPWR U$$2245/X sky130_fd_sc_hd__xor2_1
XFILLER_16_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1500 U$$950/B1 U$$1504/A2 U$$2324/A1 U$$1504/B2 VGND VGND VPWR VPWR U$$1501/A
+ sky130_fd_sc_hd__a22o_1
XU$$1511 U$$1509/Y input15/X input14/X U$$1510/X U$$1507/Y VGND VGND VPWR VPWR U$$1511/X
+ sky130_fd_sc_hd__a32o_2
XU$$2256 U$$3213/B1 U$$2302/A2 U$$477/A1 U$$2302/B2 VGND VGND VPWR VPWR U$$2257/A
+ sky130_fd_sc_hd__a22o_1
XU$$2267 U$$2267/A U$$2309/B VGND VGND VPWR VPWR U$$2267/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1522 U$$1522/A U$$1546/B VGND VGND VPWR VPWR U$$1522/X sky130_fd_sc_hd__xor2_1
XFILLER_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2278 U$$3235/B1 U$$2316/A2 U$$2691/A1 U$$2316/B2 VGND VGND VPWR VPWR U$$2279/A
+ sky130_fd_sc_hd__a22o_1
XU$$1533 U$$985/A1 U$$1545/A2 U$$987/A1 U$$1545/B2 VGND VGND VPWR VPWR U$$1534/A sky130_fd_sc_hd__a22o_1
XFILLER_62_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1544 U$$1544/A U$$1546/B VGND VGND VPWR VPWR U$$1544/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2289 U$$2289/A U$$2328/A VGND VGND VPWR VPWR U$$2289/X sky130_fd_sc_hd__xor2_1
XFILLER_43_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1555 U$$594/B1 U$$1557/A2 U$$461/A1 U$$1557/B2 VGND VGND VPWR VPWR U$$1556/A sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_116_0 dadda_ha_3_116_0/A U$$3697/X VGND VGND VPWR VPWR dadda_fa_4_117_2/CIN
+ dadda_ha_3_116_0/SUM sky130_fd_sc_hd__ha_1
XU$$1566 U$$1566/A U$$1592/B VGND VGND VPWR VPWR U$$1566/X sky130_fd_sc_hd__xor2_1
XFILLER_176_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1577 U$$1714/A1 U$$1621/A2 U$$2949/A1 U$$1621/B2 VGND VGND VPWR VPWR U$$1578/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1588 U$$1588/A U$$1620/B VGND VGND VPWR VPWR U$$1588/X sky130_fd_sc_hd__xor2_1
XFILLER_187_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1599 U$$3243/A1 U$$1607/A2 U$$3108/A1 U$$1607/B2 VGND VGND VPWR VPWR U$$1600/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_115_0 dadda_fa_7_115_0/A dadda_fa_7_115_0/B dadda_fa_7_115_0/CIN VGND
+ VGND VPWR VPWR _412_/D _283_/D sky130_fd_sc_hd__fa_1
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1014 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_60_0 dadda_fa_2_60_0/A dadda_fa_2_60_0/B dadda_fa_2_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_0/B dadda_fa_3_60_2/B sky130_fd_sc_hd__fa_1
Xrepeater400 U$$783/A2 VGND VGND VPWR VPWR U$$711/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$207 final_adder.U$$206/B final_adder.U$$977/B1 final_adder.U$$207/B1
+ VGND VGND VPWR VPWR final_adder.U$$207/X sky130_fd_sc_hd__a21o_1
XFILLER_131_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater411 U$$678/A2 VGND VGND VPWR VPWR U$$652/A2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$218 final_adder.U$$218/A final_adder.U$$218/B VGND VGND VPWR VPWR
+ final_adder.U$$346/B sky130_fd_sc_hd__and2_1
Xrepeater422 U$$4251/X VGND VGND VPWR VPWR U$$4373/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$229 final_adder.U$$228/B final_adder.U$$999/B1 final_adder.U$$229/B1
+ VGND VGND VPWR VPWR final_adder.U$$229/X sky130_fd_sc_hd__a21o_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater433 U$$4114/X VGND VGND VPWR VPWR U$$4176/A2 sky130_fd_sc_hd__buf_4
XFILLER_27_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater444 U$$134/A2 VGND VGND VPWR VPWR U$$122/A2 sky130_fd_sc_hd__buf_8
XFILLER_84_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater455 U$$3874/A2 VGND VGND VPWR VPWR U$$3878/A2 sky130_fd_sc_hd__buf_6
Xrepeater466 U$$3833/A2 VGND VGND VPWR VPWR U$$3819/A2 sky130_fd_sc_hd__buf_6
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater477 U$$3566/X VGND VGND VPWR VPWR U$$3644/A2 sky130_fd_sc_hd__buf_6
XU$$4170 U$$4307/A1 U$$4176/A2 U$$4309/A1 U$$4176/B2 VGND VGND VPWR VPWR U$$4171/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater488 U$$3348/A2 VGND VGND VPWR VPWR U$$3320/A2 sky130_fd_sc_hd__buf_4
XU$$4181 U$$4181/A U$$4239/B VGND VGND VPWR VPWR U$$4181/X sky130_fd_sc_hd__xor2_1
XFILLER_81_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater499 U$$3229/A2 VGND VGND VPWR VPWR U$$3187/A2 sky130_fd_sc_hd__buf_6
XU$$4192 U$$4466/A1 U$$4210/A2 U$$4466/B1 U$$4210/B2 VGND VGND VPWR VPWR U$$4193/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1026 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3480 U$$3480/A U$$3480/B VGND VGND VPWR VPWR U$$3480/X sky130_fd_sc_hd__xor2_1
XFILLER_207_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3491 U$$4311/B1 U$$3517/A2 U$$4176/B1 U$$3517/B2 VGND VGND VPWR VPWR U$$3492/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2790 U$$2925/B1 U$$2790/A2 U$$463/A1 U$$2790/B2 VGND VGND VPWR VPWR U$$2791/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_82_1 dadda_fa_4_82_1/A dadda_fa_4_82_1/B dadda_fa_4_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/B dadda_fa_5_82_1/B sky130_fd_sc_hd__fa_1
XFILLER_136_1008 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_75_0 dadda_fa_4_75_0/A dadda_fa_4_75_0/B dadda_fa_4_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/A dadda_fa_5_75_1/A sky130_fd_sc_hd__fa_1
XFILLER_150_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput203 c[51] VGND VGND VPWR VPWR input203/X sky130_fd_sc_hd__clkbuf_4
Xinput214 c[61] VGND VGND VPWR VPWR input214/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput225 c[71] VGND VGND VPWR VPWR input225/X sky130_fd_sc_hd__clkbuf_2
XTAP_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput236 c[81] VGND VGND VPWR VPWR input236/X sky130_fd_sc_hd__clkbuf_4
XTAP_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput247 c[91] VGND VGND VPWR VPWR input247/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$741 final_adder.U$$740/B final_adder.U$$661/X final_adder.U$$629/X
+ VGND VGND VPWR VPWR final_adder.U$$741/X sky130_fd_sc_hd__a21o_1
XTAP_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$752 final_adder.U$$784/B final_adder.U$$752/B VGND VGND VPWR VPWR
+ final_adder.U$$752/X sky130_fd_sc_hd__and2_1
XTAP_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$763 final_adder.U$$762/B final_adder.U$$683/X final_adder.U$$651/X
+ VGND VGND VPWR VPWR final_adder.U$$763/X sky130_fd_sc_hd__a21o_1
XTAP_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$602 U$$52/B1 U$$636/A2 U$$56/A1 U$$636/B2 VGND VGND VPWR VPWR U$$603/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$774 final_adder.U$$774/A final_adder.U$$774/B VGND VGND VPWR VPWR
+ final_adder.U$$774/X sky130_fd_sc_hd__and2_1
XU$$613 U$$613/A U$$617/B VGND VGND VPWR VPWR U$$613/X sky130_fd_sc_hd__xor2_1
XFILLER_57_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$785 final_adder.U$$784/B final_adder.U$$705/X final_adder.U$$673/X
+ VGND VGND VPWR VPWR final_adder.U$$785/X sky130_fd_sc_hd__a21o_1
XU$$624 U$$759/B1 U$$624/A2 U$$763/A1 U$$624/B2 VGND VGND VPWR VPWR U$$625/A sky130_fd_sc_hd__a22o_1
XFILLER_44_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$796 final_adder.U$$796/A final_adder.U$$796/B VGND VGND VPWR VPWR
+ final_adder.U$$796/X sky130_fd_sc_hd__and2_1
XFILLER_44_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$635 U$$635/A U$$637/B VGND VGND VPWR VPWR U$$635/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$646 U$$920/A1 U$$652/A2 U$$783/B1 U$$652/B2 VGND VGND VPWR VPWR U$$647/A sky130_fd_sc_hd__a22o_1
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$657 U$$657/A U$$684/A VGND VGND VPWR VPWR U$$657/X sky130_fd_sc_hd__xor2_1
XFILLER_189_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$668 U$$940/B1 U$$672/A2 U$$807/A1 U$$668/B2 VGND VGND VPWR VPWR U$$669/A sky130_fd_sc_hd__a22o_1
XU$$679 U$$679/A U$$684/A VGND VGND VPWR VPWR U$$679/X sky130_fd_sc_hd__xor2_1
XFILLER_44_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1502 U$$4103/B1 VGND VGND VPWR VPWR U$$4379/A1 sky130_fd_sc_hd__buf_6
Xrepeater1513 U$$950/A1 VGND VGND VPWR VPWR U$$676/A1 sky130_fd_sc_hd__buf_4
XFILLER_197_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1524 U$$3578/B1 VGND VGND VPWR VPWR U$$3032/A1 sky130_fd_sc_hd__buf_4
Xrepeater1535 U$$3/A VGND VGND VPWR VPWR U$$127/B sky130_fd_sc_hd__buf_6
Xrepeater1546 U$$3684/B1 VGND VGND VPWR VPWR U$$3547/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1557 U$$1764/B1 VGND VGND VPWR VPWR U$$944/A1 sky130_fd_sc_hd__buf_6
XFILLER_99_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1568 U$$4504/A1 VGND VGND VPWR VPWR U$$2449/A1 sky130_fd_sc_hd__buf_6
Xrepeater1579 U$$116/A1 VGND VGND VPWR VPWR U$$388/B1 sky130_fd_sc_hd__buf_8
XFILLER_153_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2020 U$$787/A1 U$$2052/A2 U$$652/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2021/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_32_4 U$$1667/X U$$1800/X U$$1933/X VGND VGND VPWR VPWR dadda_fa_3_33_1/CIN
+ dadda_fa_3_32_3/CIN sky130_fd_sc_hd__fa_1
XU$$2031 U$$2031/A U$$2047/B VGND VGND VPWR VPWR U$$2031/X sky130_fd_sc_hd__xor2_1
XU$$2042 U$$4508/A1 U$$1922/X U$$948/A1 U$$1923/X VGND VGND VPWR VPWR U$$2043/A sky130_fd_sc_hd__a22o_1
XFILLER_165_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2053 U$$2053/A U$$2054/A VGND VGND VPWR VPWR U$$2053/X sky130_fd_sc_hd__xor2_1
XFILLER_23_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2064 U$$2064/A U$$2094/B VGND VGND VPWR VPWR U$$2064/X sky130_fd_sc_hd__xor2_1
XFILLER_200_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1330 U$$1330/A U$$1330/B VGND VGND VPWR VPWR U$$1330/X sky130_fd_sc_hd__xor2_1
XU$$2075 U$$3719/A1 U$$2093/A2 U$$3447/A1 U$$2093/B2 VGND VGND VPWR VPWR U$$2076/A
+ sky130_fd_sc_hd__a22o_1
XU$$2086 U$$2086/A U$$2092/B VGND VGND VPWR VPWR U$$2086/X sky130_fd_sc_hd__xor2_1
XU$$1341 U$$2026/A1 U$$1353/A2 U$$932/A1 U$$1349/B2 VGND VGND VPWR VPWR U$$1342/A
+ sky130_fd_sc_hd__a22o_1
XU$$2097 U$$4289/A1 U$$2099/A2 U$$3878/B1 U$$2099/B2 VGND VGND VPWR VPWR U$$2098/A
+ sky130_fd_sc_hd__a22o_1
XU$$1352 U$$1352/A U$$1366/B VGND VGND VPWR VPWR U$$1352/X sky130_fd_sc_hd__xor2_1
XFILLER_210_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1363 U$$950/B1 U$$1367/A2 U$$2324/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1364/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1374 U$$1372/Y input13/X U$$1370/A U$$1373/X U$$1370/Y VGND VGND VPWR VPWR U$$1374/X
+ sky130_fd_sc_hd__a32o_4
XU$$1385 U$$1385/A U$$1399/B VGND VGND VPWR VPWR U$$1385/X sky130_fd_sc_hd__xor2_1
XFILLER_149_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1396 U$$985/A1 U$$1404/A2 U$$987/A1 U$$1404/B2 VGND VGND VPWR VPWR U$$1397/A sky130_fd_sc_hd__a22o_1
XFILLER_149_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_92_0 dadda_fa_5_92_0/A dadda_fa_5_92_0/B dadda_fa_5_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_93_0/A dadda_fa_6_92_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_209_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_77_6 U$$3752/X U$$3885/X U$$4018/X VGND VGND VPWR VPWR dadda_fa_2_78_2/B
+ dadda_fa_2_77_5/B sky130_fd_sc_hd__fa_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_353 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_887 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$70 _366_/Q _238_/Q VGND VGND VPWR VPWR final_adder.U$$955/B1 final_adder.U$$184/A
+ sky130_fd_sc_hd__ha_1
XFILLER_14_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$81 _377_/Q _249_/Q VGND VGND VPWR VPWR final_adder.U$$175/B1 final_adder.U$$174/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$92 _388_/Q _260_/Q VGND VGND VPWR VPWR final_adder.U$$933/B1 final_adder.U$$162/A
+ sky130_fd_sc_hd__ha_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_439 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_101_1 input131/X dadda_fa_3_101_1/B dadda_fa_3_101_1/CIN VGND VGND VPWR
+ VPWR dadda_fa_4_102_0/CIN dadda_fa_4_101_2/A sky130_fd_sc_hd__fa_1
XFILLER_102_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_118_0_1868 VGND VGND VPWR VPWR dadda_fa_4_118_0/A dadda_fa_4_118_0_1868/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_27_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_122_0 dadda_fa_6_122_0/A dadda_fa_6_122_0/B dadda_fa_6_122_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_123_0/B dadda_fa_7_122_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_65_4 U$$1733/X U$$1866/X U$$1999/X VGND VGND VPWR VPWR dadda_fa_1_66_6/CIN
+ dadda_fa_1_65_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_42_3 dadda_fa_3_42_3/A dadda_fa_3_42_3/B dadda_fa_3_42_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_43_1/B dadda_fa_4_42_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_36_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$560 final_adder.U$$568/B final_adder.U$$560/B VGND VGND VPWR VPWR
+ final_adder.U$$680/B sky130_fd_sc_hd__and2_1
XFILLER_188_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$571 final_adder.U$$570/B final_adder.U$$455/X final_adder.U$$447/X
+ VGND VGND VPWR VPWR final_adder.U$$571/X sky130_fd_sc_hd__a21o_1
XTAP_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$410 U$$410/A VGND VGND VPWR VPWR U$$410/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$582 final_adder.U$$590/B final_adder.U$$582/B VGND VGND VPWR VPWR
+ final_adder.U$$702/B sky130_fd_sc_hd__and2_1
XTAP_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$421 U$$8/B1 U$$437/A2 U$$12/A1 U$$437/B2 VGND VGND VPWR VPWR U$$422/A sky130_fd_sc_hd__a22o_1
XTAP_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_35_2 dadda_fa_3_35_2/A dadda_fa_3_35_2/B dadda_fa_3_35_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_1/A dadda_fa_4_35_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$593 final_adder.U$$592/B final_adder.U$$477/X final_adder.U$$469/X
+ VGND VGND VPWR VPWR final_adder.U$$593/X sky130_fd_sc_hd__a21o_1
XU$$432 U$$432/A U$$516/B VGND VGND VPWR VPWR U$$432/X sky130_fd_sc_hd__xor2_1
XTAP_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$443 U$$717/A1 U$$515/A2 U$$34/A1 U$$515/B2 VGND VGND VPWR VPWR U$$444/A sky130_fd_sc_hd__a22o_1
XTAP_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$454 U$$454/A U$$474/B VGND VGND VPWR VPWR U$$454/X sky130_fd_sc_hd__xor2_1
XFILLER_189_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_28_1 U$$1925/X U$$1993/B input177/X VGND VGND VPWR VPWR dadda_fa_4_29_0/CIN
+ dadda_fa_4_28_2/A sky130_fd_sc_hd__fa_1
XFILLER_17_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$465 U$$54/A1 U$$483/A2 U$$56/A1 U$$483/B2 VGND VGND VPWR VPWR U$$466/A sky130_fd_sc_hd__a22o_1
XFILLER_205_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$476 U$$476/A U$$504/B VGND VGND VPWR VPWR U$$476/X sky130_fd_sc_hd__xor2_1
XU$$487 U$$759/B1 U$$491/A2 U$$763/A1 U$$491/B2 VGND VGND VPWR VPWR U$$488/A sky130_fd_sc_hd__a22o_1
XU$$498 U$$498/A U$$536/B VGND VGND VPWR VPWR U$$498/X sky130_fd_sc_hd__xor2_1
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_970 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1310 U$$3377/B VGND VGND VPWR VPWR U$$3375/B sky130_fd_sc_hd__buf_8
Xrepeater1321 input42/X VGND VGND VPWR VPWR U$$3288/A sky130_fd_sc_hd__buf_4
XFILLER_5_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1332 U$$2950/B VGND VGND VPWR VPWR U$$2920/B sky130_fd_sc_hd__buf_8
XFILLER_125_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1343 U$$2837/B VGND VGND VPWR VPWR U$$2825/B sky130_fd_sc_hd__buf_6
XFILLER_125_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1354 U$$260/B VGND VGND VPWR VPWR U$$244/B sky130_fd_sc_hd__buf_8
XFILLER_153_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_87_5 dadda_fa_2_87_5/A dadda_fa_2_87_5/B dadda_fa_2_87_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_88_2/A dadda_fa_4_87_0/A sky130_fd_sc_hd__fa_1
Xrepeater1365 input33/X VGND VGND VPWR VPWR U$$2716/B sky130_fd_sc_hd__buf_8
XFILLER_126_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1376 U$$794/B VGND VGND VPWR VPWR U$$784/B sky130_fd_sc_hd__buf_6
Xrepeater1387 U$$2466/A VGND VGND VPWR VPWR U$$2442/B sky130_fd_sc_hd__buf_6
XFILLER_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1398 input27/X VGND VGND VPWR VPWR U$$2317/B sky130_fd_sc_hd__buf_8
XFILLER_80_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_30_1 U$$466/X U$$599/X U$$732/X VGND VGND VPWR VPWR dadda_fa_3_31_1/B
+ dadda_fa_3_30_3/A sky130_fd_sc_hd__fa_1
XFILLER_51_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1160 U$$62/B1 U$$1204/A2 U$$888/A1 U$$1204/B2 VGND VGND VPWR VPWR U$$1161/A sky130_fd_sc_hd__a22o_1
XU$$1171 U$$1171/A U$$1175/B VGND VGND VPWR VPWR U$$1171/X sky130_fd_sc_hd__xor2_1
XU$$1182 U$$3922/A1 U$$1222/A2 U$$3922/B1 U$$1222/B2 VGND VGND VPWR VPWR U$$1183/A
+ sky130_fd_sc_hd__a22o_1
XU$$1193 U$$1193/A U$$1205/B VGND VGND VPWR VPWR U$$1193/X sky130_fd_sc_hd__xor2_1
XFILLER_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_117_1 dadda_fa_5_117_1/A dadda_fa_5_117_1/B dadda_fa_5_117_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_118_0/B dadda_fa_7_117_0/A sky130_fd_sc_hd__fa_1
XFILLER_108_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1092 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_82_4 U$$2831/X U$$2964/X U$$3097/X VGND VGND VPWR VPWR dadda_fa_2_83_2/CIN
+ dadda_fa_2_82_5/A sky130_fd_sc_hd__fa_1
XFILLER_104_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_75_3 U$$2817/X U$$2950/X U$$3083/X VGND VGND VPWR VPWR dadda_fa_2_76_1/B
+ dadda_fa_2_75_4/B sky130_fd_sc_hd__fa_1
XFILLER_120_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_52_2 dadda_fa_4_52_2/A dadda_fa_4_52_2/B dadda_fa_4_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_53_0/CIN dadda_fa_5_52_1/CIN sky130_fd_sc_hd__fa_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_2 U$$3335/X U$$3468/X U$$3601/X VGND VGND VPWR VPWR dadda_fa_2_69_1/A
+ dadda_fa_2_68_4/A sky130_fd_sc_hd__fa_1
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_45_1 dadda_fa_4_45_1/A dadda_fa_4_45_1/B dadda_fa_4_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/B dadda_fa_5_45_1/B sky130_fd_sc_hd__fa_1
XFILLER_65_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_22_0 dadda_fa_7_22_0/A dadda_fa_7_22_0/B dadda_fa_7_22_0/CIN VGND VGND
+ VPWR VPWR _319_/D _190_/D sky130_fd_sc_hd__fa_2
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_38_0 dadda_fa_4_38_0/A dadda_fa_4_38_0/B dadda_fa_4_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/A dadda_fa_5_38_1/A sky130_fd_sc_hd__fa_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _384_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _420_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 input254/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 U$$3207/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _351_/CLK _350_/D VGND VGND VPWR VPWR _350_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_281_ _411_/CLK _281_/D VGND VGND VPWR VPWR _281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_57_2 U$$919/X U$$1052/X VGND VGND VPWR VPWR dadda_fa_1_58_7/CIN dadda_fa_2_57_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_190_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_70_2 U$$1211/X U$$1344/X U$$1477/X VGND VGND VPWR VPWR dadda_fa_1_71_7/A
+ dadda_fa_1_70_8/B sky130_fd_sc_hd__fa_1
XTAP_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_754 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_1 U$$532/X U$$665/X U$$798/X VGND VGND VPWR VPWR dadda_fa_1_64_5/CIN
+ dadda_fa_1_63_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_37_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_40_0 dadda_fa_3_40_0/A dadda_fa_3_40_0/B dadda_fa_3_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_0/B dadda_fa_4_40_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_56_0 U$$119/X U$$252/X U$$385/X VGND VGND VPWR VPWR dadda_fa_1_57_7/B
+ dadda_fa_1_56_8/B sky130_fd_sc_hd__fa_1
XTAP_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$390 final_adder.U$$394/B final_adder.U$$390/B VGND VGND VPWR VPWR
+ final_adder.U$$514/B sky130_fd_sc_hd__and2_2
XFILLER_188_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$240 U$$240/A U$$244/B VGND VGND VPWR VPWR U$$240/X sky130_fd_sc_hd__xor2_1
XFILLER_206_955 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$251 U$$251/A1 U$$257/A2 U$$388/B1 U$$257/B2 VGND VGND VPWR VPWR U$$252/A sky130_fd_sc_hd__a22o_1
XFILLER_45_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$262 U$$262/A U$$272/B VGND VGND VPWR VPWR U$$262/X sky130_fd_sc_hd__xor2_1
XFILLER_73_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$273 U$$274/A VGND VGND VPWR VPWR U$$273/Y sky130_fd_sc_hd__inv_1
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$284 U$$8/B1 U$$316/A2 U$$12/A1 U$$316/B2 VGND VGND VPWR VPWR U$$285/A sky130_fd_sc_hd__a22o_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$295 U$$295/A U$$379/B VGND VGND VPWR VPWR U$$295/X sky130_fd_sc_hd__xor2_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1 U$$1/A VGND VGND VPWR VPWR U$$3/B sky130_fd_sc_hd__inv_1
XFILLER_199_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$9 _305_/Q _177_/Q VGND VGND VPWR VPWR final_adder.U$$9/COUT final_adder.U$$9/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_65_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput304 output304/A VGND VGND VPWR VPWR o[27] sky130_fd_sc_hd__buf_2
XFILLER_161_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_92_3 U$$4181/X U$$4314/X U$$4447/X VGND VGND VPWR VPWR dadda_fa_3_93_1/B
+ dadda_fa_3_92_3/B sky130_fd_sc_hd__fa_1
Xoutput315 output315/A VGND VGND VPWR VPWR o[37] sky130_fd_sc_hd__buf_2
XFILLER_99_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput326 output326/A VGND VGND VPWR VPWR o[47] sky130_fd_sc_hd__buf_2
Xrepeater1140 U$$721/B1 VGND VGND VPWR VPWR U$$997/A1 sky130_fd_sc_hd__buf_6
XFILLER_99_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput337 output337/A VGND VGND VPWR VPWR o[57] sky130_fd_sc_hd__buf_2
XFILLER_142_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1151 U$$4144/B1 VGND VGND VPWR VPWR U$$4420/A1 sky130_fd_sc_hd__buf_8
Xrepeater1162 input7/X VGND VGND VPWR VPWR U$$962/A sky130_fd_sc_hd__buf_4
Xdadda_fa_2_85_2 dadda_fa_2_85_2/A dadda_fa_2_85_2/B dadda_fa_2_85_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/A dadda_fa_3_85_3/A sky130_fd_sc_hd__fa_1
Xoutput348 output348/A VGND VGND VPWR VPWR o[67] sky130_fd_sc_hd__buf_2
XFILLER_82_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput359 output359/A VGND VGND VPWR VPWR o[77] sky130_fd_sc_hd__buf_2
XFILLER_142_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1173 U$$3183/A1 VGND VGND VPWR VPWR U$$991/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1184 input67/X VGND VGND VPWR VPWR U$$30/A1 sky130_fd_sc_hd__buf_4
XFILLER_142_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_62_1 dadda_fa_5_62_1/A dadda_fa_5_62_1/B dadda_fa_5_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_63_0/B dadda_fa_7_62_0/A sky130_fd_sc_hd__fa_2
Xrepeater1195 U$$4410/B1 VGND VGND VPWR VPWR U$$4275/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_78_1 dadda_fa_2_78_1/A dadda_fa_2_78_1/B dadda_fa_2_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_0/CIN dadda_fa_3_78_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_55_0 dadda_fa_5_55_0/A dadda_fa_5_55_0/B dadda_fa_5_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_56_0/A dadda_fa_6_55_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_45_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_54_8 input206/X dadda_fa_1_54_8/B dadda_fa_1_54_8/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_55_3/A dadda_fa_3_54_0/A sky130_fd_sc_hd__fa_2
XFILLER_56_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_101_0 U$$2602/Y U$$2736/X U$$2869/X VGND VGND VPWR VPWR dadda_fa_3_102_1/CIN
+ dadda_fa_3_101_3/A sky130_fd_sc_hd__fa_1
XFILLER_63_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_80_1 U$$1497/X U$$1630/X U$$1763/X VGND VGND VPWR VPWR dadda_fa_2_81_1/A
+ dadda_fa_2_80_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_73_0 U$$1882/X U$$2015/X U$$2148/X VGND VGND VPWR VPWR dadda_fa_2_74_0/B
+ dadda_fa_2_73_3/B sky130_fd_sc_hd__fa_1
XFILLER_28_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3309 U$$3309/A U$$3395/B VGND VGND VPWR VPWR U$$3309/X sky130_fd_sc_hd__xor2_1
XFILLER_86_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2608 U$$2606/B input31/X input32/X U$$2603/Y VGND VGND VPWR VPWR U$$2608/X sky130_fd_sc_hd__a22o_4
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_640 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2619 U$$2754/B1 U$$2625/A2 U$$2621/A1 U$$2625/B2 VGND VGND VPWR VPWR U$$2620/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1907 U$$948/A1 U$$1785/X U$$2044/B1 U$$1786/X VGND VGND VPWR VPWR U$$1908/A sky130_fd_sc_hd__a22o_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1918 input20/X VGND VGND VPWR VPWR U$$1918/Y sky130_fd_sc_hd__inv_1
XFILLER_54_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ _408_/CLK _402_/D VGND VGND VPWR VPWR _402_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1929 U$$1929/A U$$1991/B VGND VGND VPWR VPWR U$$1929/X sky130_fd_sc_hd__xor2_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_333_ _342_/CLK _333_/D VGND VGND VPWR VPWR _333_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_264_ _401_/CLK _264_/D VGND VGND VPWR VPWR _264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_195_ _323_/CLK _195_/D VGND VGND VPWR VPWR _195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_95_1 dadda_fa_3_95_1/A dadda_fa_3_95_1/B dadda_fa_3_95_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_0/CIN dadda_fa_4_95_2/A sky130_fd_sc_hd__fa_1
XFILLER_143_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_72_0 dadda_fa_6_72_0/A dadda_fa_6_72_0/B dadda_fa_6_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_73_0/B dadda_fa_7_72_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_88_0 dadda_fa_3_88_0/A dadda_fa_3_88_0/B dadda_fa_3_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_0/B dadda_fa_4_88_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_9_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater807 U$$2252/B2 VGND VGND VPWR VPWR U$$2226/B2 sky130_fd_sc_hd__buf_6
Xrepeater818 U$$2169/B2 VGND VGND VPWR VPWR U$$2149/B2 sky130_fd_sc_hd__buf_6
XU$$4500 U$$4500/A1 U$$4388/X U$$4502/A1 U$$4512/B2 VGND VGND VPWR VPWR U$$4501/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater829 U$$1923/X VGND VGND VPWR VPWR U$$2040/B2 sky130_fd_sc_hd__buf_4
XFILLER_42_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4511 U$$4511/A U$$4511/B VGND VGND VPWR VPWR U$$4511/X sky130_fd_sc_hd__xor2_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$14 U$$14/A1 U$$8/A2 U$$16/A1 U$$8/B2 VGND VGND VPWR VPWR U$$15/A sky130_fd_sc_hd__a22o_1
XU$$3810 U$$3810/A U$$3814/B VGND VGND VPWR VPWR U$$3810/X sky130_fd_sc_hd__xor2_1
XU$$25 U$$25/A U$$9/B VGND VGND VPWR VPWR U$$25/X sky130_fd_sc_hd__xor2_1
XU$$3821 input117/X U$$3833/A2 input118/X U$$3833/B2 VGND VGND VPWR VPWR U$$3822/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_117_0 U$$3698/Y U$$3832/X U$$3965/X VGND VGND VPWR VPWR dadda_fa_5_118_0/A
+ dadda_fa_5_117_1/A sky130_fd_sc_hd__fa_1
XTAP_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$36 U$$36/A1 U$$42/A2 U$$38/A1 U$$42/B2 VGND VGND VPWR VPWR U$$37/A sky130_fd_sc_hd__a22o_1
XU$$3832 U$$3832/A U$$3834/B VGND VGND VPWR VPWR U$$3832/X sky130_fd_sc_hd__xor2_1
XTAP_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$47 U$$47/A U$$51/B VGND VGND VPWR VPWR U$$47/X sky130_fd_sc_hd__xor2_1
XTAP_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3843 U$$3843/A U$$3927/B VGND VGND VPWR VPWR U$$3843/X sky130_fd_sc_hd__xor2_1
XU$$58 U$$58/A1 U$$94/A2 U$$60/A1 U$$94/B2 VGND VGND VPWR VPWR U$$59/A sky130_fd_sc_hd__a22o_1
XU$$3854 U$$4402/A1 U$$3874/A2 U$$4402/B1 U$$3874/B2 VGND VGND VPWR VPWR U$$3855/A
+ sky130_fd_sc_hd__a22o_1
XU$$69 U$$69/A U$$81/B VGND VGND VPWR VPWR U$$69/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_5_4_0 U$$15/X U$$148/X VGND VGND VPWR VPWR dadda_fa_6_5_0/CIN dadda_fa_7_4_0/A
+ sky130_fd_sc_hd__ha_1
XU$$3865 U$$3865/A U$$3903/B VGND VGND VPWR VPWR U$$3865/X sky130_fd_sc_hd__xor2_1
XFILLER_24_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3876 U$$4424/A1 U$$3878/A2 U$$3876/B1 U$$3878/B2 VGND VGND VPWR VPWR U$$3877/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3887 U$$3887/A U$$3971/B VGND VGND VPWR VPWR U$$3887/X sky130_fd_sc_hd__xor2_1
XTAP_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3898 U$$4309/A1 U$$3902/A2 U$$4309/B1 U$$3902/B2 VGND VGND VPWR VPWR U$$3899/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4503_1828 VGND VGND VPWR VPWR U$$4503_1828/HI U$$4503/B sky130_fd_sc_hd__conb_1
XFILLER_21_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_16 _328_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_27 _337_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_38 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 _341_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_832 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_898 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4395_1774 VGND VGND VPWR VPWR U$$4395_1774/HI U$$4395/B sky130_fd_sc_hd__conb_1
Xdadda_fa_2_90_0 U$$3246/X U$$3379/X U$$3512/X VGND VGND VPWR VPWR dadda_fa_3_91_0/B
+ dadda_fa_3_90_2/B sky130_fd_sc_hd__fa_1
XFILLER_127_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_46_6 U$$2493/X U$$2626/X VGND VGND VPWR VPWR dadda_fa_2_47_3/CIN dadda_fa_3_46_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_114_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_52_5 U$$2372/X U$$2505/X U$$2638/X VGND VGND VPWR VPWR dadda_fa_2_53_2/A
+ dadda_fa_2_52_5/A sky130_fd_sc_hd__fa_1
XFILLER_110_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_45_4 U$$1693/X U$$1826/X U$$1959/X VGND VGND VPWR VPWR dadda_fa_2_46_3/B
+ dadda_fa_2_45_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_15_2 input163/X dadda_fa_4_15_2/B dadda_ha_3_15_0/SUM VGND VGND VPWR VPWR
+ dadda_fa_5_16_0/CIN dadda_fa_5_15_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$1019 final_adder.U$$6/SUM final_adder.U$$505/X final_adder.U$$6/COUT
+ VGND VGND VPWR VPWR final_adder.U$$1031/B sky130_fd_sc_hd__a21o_1
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3106 U$$3243/A1 U$$3108/A2 U$$3108/A1 U$$3108/B2 VGND VGND VPWR VPWR U$$3107/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_1140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3117 U$$3117/A U$$3117/B VGND VGND VPWR VPWR U$$3117/X sky130_fd_sc_hd__xor2_1
XFILLER_47_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3128 U$$251/A1 U$$3132/A2 U$$116/A1 U$$3132/B2 VGND VGND VPWR VPWR U$$3129/A sky130_fd_sc_hd__a22o_1
XU$$3139 U$$3139/A U$$3150/A VGND VGND VPWR VPWR U$$3139/X sky130_fd_sc_hd__xor2_1
XFILLER_100_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2405 U$$896/B1 U$$2435/A2 U$$3366/A1 U$$2435/B2 VGND VGND VPWR VPWR U$$2406/A
+ sky130_fd_sc_hd__a22o_1
XU$$2416 U$$2416/A U$$2426/B VGND VGND VPWR VPWR U$$2416/X sky130_fd_sc_hd__xor2_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2427 U$$3112/A1 U$$2449/A2 U$$3114/A1 U$$2449/B2 VGND VGND VPWR VPWR U$$2428/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2438 U$$2438/A U$$2442/B VGND VGND VPWR VPWR U$$2438/X sky130_fd_sc_hd__xor2_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1704 U$$2113/B1 U$$1706/A2 U$$3348/B1 U$$1706/B2 VGND VGND VPWR VPWR U$$1705/A
+ sky130_fd_sc_hd__a22o_1
XU$$2449 U$$2449/A1 U$$2449/A2 U$$4506/A1 U$$2449/B2 VGND VGND VPWR VPWR U$$2450/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1715 U$$1715/A U$$1721/B VGND VGND VPWR VPWR U$$1715/X sky130_fd_sc_hd__xor2_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1726 U$$630/A1 U$$1736/A2 U$$630/B1 U$$1736/B2 VGND VGND VPWR VPWR U$$1727/A sky130_fd_sc_hd__a22o_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1737 U$$1737/A U$$1739/B VGND VGND VPWR VPWR U$$1737/X sky130_fd_sc_hd__xor2_1
XFILLER_14_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1748 U$$789/A1 U$$1764/A2 U$$928/A1 U$$1764/B2 VGND VGND VPWR VPWR U$$1749/A sky130_fd_sc_hd__a22o_1
XFILLER_187_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1759 U$$1759/A U$$1765/B VGND VGND VPWR VPWR U$$1759/X sky130_fd_sc_hd__xor2_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_316_ _326_/CLK _316_/D VGND VGND VPWR VPWR _316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_247_ _377_/CLK _247_/D VGND VGND VPWR VPWR _247_/Q sky130_fd_sc_hd__dfxtp_1
Xinput14 a[21] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__buf_2
XFILLER_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput25 a[31] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__buf_6
XFILLER_155_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput36 a[41] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__buf_4
XFILLER_196_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput47 a[51] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__buf_2
Xinput58 a[61] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_178_ _327_/CLK _178_/D VGND VGND VPWR VPWR _178_/Q sky130_fd_sc_hd__dfxtp_1
Xinput69 b[13] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__buf_6
XFILLER_128_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_1166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_62_4 dadda_fa_2_62_4/A dadda_fa_2_62_4/B dadda_fa_2_62_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_1/CIN dadda_fa_3_62_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater604 U$$1591/A2 VGND VGND VPWR VPWR U$$1557/A2 sky130_fd_sc_hd__buf_6
XFILLER_81_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater615 U$$141/X VGND VGND VPWR VPWR U$$263/A2 sky130_fd_sc_hd__buf_6
XFILLER_46_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater626 U$$1353/A2 VGND VGND VPWR VPWR U$$1323/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_55_3 dadda_fa_2_55_3/A dadda_fa_2_55_3/B dadda_fa_2_55_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/B dadda_fa_3_55_3/B sky130_fd_sc_hd__fa_1
Xrepeater637 U$$1100/X VGND VGND VPWR VPWR U$$1230/A2 sky130_fd_sc_hd__buf_6
XFILLER_78_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4330 U$$4330/A U$$4330/B VGND VGND VPWR VPWR U$$4330/X sky130_fd_sc_hd__xor2_1
Xrepeater648 U$$882/B2 VGND VGND VPWR VPWR U$$872/B2 sky130_fd_sc_hd__clkbuf_4
XU$$4341 U$$4478/A1 U$$4349/A2 U$$4478/B1 U$$4349/B2 VGND VGND VPWR VPWR U$$4342/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater659 U$$759/B2 VGND VGND VPWR VPWR U$$749/B2 sky130_fd_sc_hd__buf_6
XFILLER_38_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4352 U$$4352/A input60/X VGND VGND VPWR VPWR U$$4352/X sky130_fd_sc_hd__xor2_1
XFILLER_42_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_48_2 dadda_fa_2_48_2/A dadda_fa_2_48_2/B dadda_fa_2_48_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/A dadda_fa_3_48_3/A sky130_fd_sc_hd__fa_1
XU$$4363 U$$4500/A1 U$$4373/A2 U$$4502/A1 U$$4373/B2 VGND VGND VPWR VPWR U$$4364/A
+ sky130_fd_sc_hd__a22o_1
XU$$4374 U$$4374/A input60/X VGND VGND VPWR VPWR U$$4374/X sky130_fd_sc_hd__xor2_1
XFILLER_203_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4385 U$$4385/A VGND VGND VPWR VPWR U$$4387/B sky130_fd_sc_hd__inv_1
XU$$3640 U$$3775/B1 U$$3566/X U$$3642/A1 U$$3567/X VGND VGND VPWR VPWR U$$3641/A sky130_fd_sc_hd__a22o_1
XU$$3651 U$$3651/A U$$3683/B VGND VGND VPWR VPWR U$$3651/X sky130_fd_sc_hd__xor2_1
XU$$4396 U$$4396/A1 U$$4388/X U$$4398/A1 U$$4432/B2 VGND VGND VPWR VPWR U$$4397/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_25_1 dadda_fa_5_25_1/A dadda_fa_5_25_1/B dadda_fa_5_25_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_26_0/B dadda_fa_7_25_0/A sky130_fd_sc_hd__fa_2
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3662 U$$4210/A1 U$$3680/A2 U$$4210/B1 U$$3680/B2 VGND VGND VPWR VPWR U$$3663/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3673 U$$3673/A U$$3683/B VGND VGND VPWR VPWR U$$3673/X sky130_fd_sc_hd__xor2_1
XU$$3684 U$$3684/A1 U$$3686/A2 U$$3684/B1 U$$3686/B2 VGND VGND VPWR VPWR U$$3685/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_18_0 dadda_fa_5_18_0/A dadda_fa_5_18_0/B dadda_fa_5_18_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_19_0/A dadda_fa_6_18_0/CIN sky130_fd_sc_hd__fa_1
XU$$3695 U$$3695/A U$$3698/A VGND VGND VPWR VPWR U$$3695/X sky130_fd_sc_hd__xor2_1
XU$$2950 U$$2950/A U$$2950/B VGND VGND VPWR VPWR U$$2950/X sky130_fd_sc_hd__xor2_1
XU$$2961 U$$3644/B1 U$$2985/A2 U$$3511/A1 U$$2985/B2 VGND VGND VPWR VPWR U$$2962/A
+ sky130_fd_sc_hd__a22o_1
XU$$2972 U$$2972/A U$$2978/B VGND VGND VPWR VPWR U$$2972/X sky130_fd_sc_hd__xor2_1
XU$$2983 U$$4490/A1 U$$2985/A2 U$$4492/A1 U$$2985/B2 VGND VGND VPWR VPWR U$$2984/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2994 U$$2994/A U$$2996/B VGND VGND VPWR VPWR U$$2994/X sky130_fd_sc_hd__xor2_1
XFILLER_194_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$901 final_adder.U$$130/A final_adder.U$$839/X final_adder.U$$901/B1
+ VGND VGND VPWR VPWR final_adder.U$$901/X sky130_fd_sc_hd__a21o_1
XTAP_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$923 final_adder.U$$152/A final_adder.U$$861/X final_adder.U$$923/B1
+ VGND VGND VPWR VPWR final_adder.U$$923/X sky130_fd_sc_hd__a21o_1
XFILLER_180_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$945 final_adder.U$$174/A final_adder.U$$883/X final_adder.U$$945/B1
+ VGND VGND VPWR VPWR final_adder.U$$945/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_2 U$$905/X U$$1038/X U$$1171/X VGND VGND VPWR VPWR dadda_fa_2_51_1/A
+ dadda_fa_2_50_4/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$967 final_adder.U$$196/A final_adder.U$$809/X final_adder.U$$967/B1
+ VGND VGND VPWR VPWR final_adder.U$$967/X sky130_fd_sc_hd__a21o_1
XU$$806 U$$806/A U$$808/B VGND VGND VPWR VPWR U$$806/X sky130_fd_sc_hd__xor2_1
XFILLER_56_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$817 U$$954/A1 U$$689/X U$$817/B1 U$$690/X VGND VGND VPWR VPWR U$$818/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_43_1 U$$492/X U$$625/X U$$758/X VGND VGND VPWR VPWR dadda_fa_2_44_3/A
+ dadda_fa_2_43_5/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$989 final_adder.U$$218/A final_adder.U$$831/X final_adder.U$$989/B1
+ VGND VGND VPWR VPWR final_adder.U$$989/X sky130_fd_sc_hd__a21o_1
XU$$828 U$$828/A1 U$$918/A2 U$$967/A1 U$$918/B2 VGND VGND VPWR VPWR U$$829/A sky130_fd_sc_hd__a22o_1
XFILLER_28_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$839 U$$839/A U$$847/B VGND VGND VPWR VPWR U$$839/X sky130_fd_sc_hd__xor2_1
XFILLER_84_896 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_20_0 U$$1405/B input169/X dadda_fa_4_20_0/CIN VGND VGND VPWR VPWR dadda_fa_5_21_0/A
+ dadda_fa_5_20_1/A sky130_fd_sc_hd__fa_1
XFILLER_204_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_36_0 U$$79/X U$$212/X U$$345/X VGND VGND VPWR VPWR dadda_fa_2_37_5/A dadda_fa_2_36_5/CIN
+ sky130_fd_sc_hd__fa_1
XFILLER_71_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_900 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1706 U$$4335/B1 VGND VGND VPWR VPWR U$$3378/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_153_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_72_3 dadda_fa_3_72_3/A dadda_fa_3_72_3/B dadda_fa_3_72_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_73_1/B dadda_fa_4_72_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_79_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_65_2 dadda_fa_3_65_2/A dadda_fa_3_65_2/B dadda_fa_3_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_1/A dadda_fa_4_65_2/B sky130_fd_sc_hd__fa_1
XFILLER_117_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_58_1 dadda_fa_3_58_1/A dadda_fa_3_58_1/B dadda_fa_3_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_0/CIN dadda_fa_4_58_2/A sky130_fd_sc_hd__fa_1
XFILLER_94_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_35_0 dadda_fa_6_35_0/A dadda_fa_6_35_0/B dadda_fa_6_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_36_0/B dadda_fa_7_35_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2202 U$$2202/A1 U$$2252/A2 U$$2202/B1 U$$2252/B2 VGND VGND VPWR VPWR U$$2203/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2213 U$$2213/A U$$2227/B VGND VGND VPWR VPWR U$$2213/X sky130_fd_sc_hd__xor2_1
XU$$2224 U$$3594/A1 U$$2272/A2 U$$4005/B1 U$$2272/B2 VGND VGND VPWR VPWR U$$2225/A
+ sky130_fd_sc_hd__a22o_1
XU$$2235 U$$2235/A U$$2285/B VGND VGND VPWR VPWR U$$2235/X sky130_fd_sc_hd__xor2_1
XU$$2246 U$$3614/B1 U$$2284/A2 U$$3481/A1 U$$2284/B2 VGND VGND VPWR VPWR U$$2247/A
+ sky130_fd_sc_hd__a22o_1
XU$$1501 U$$1501/A U$$1501/B VGND VGND VPWR VPWR U$$1501/X sky130_fd_sc_hd__xor2_1
XU$$1512 U$$1510/B input14/X input15/X U$$1507/Y VGND VGND VPWR VPWR U$$1512/X sky130_fd_sc_hd__a22o_2
XFILLER_16_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2257 U$$2257/A U$$2303/B VGND VGND VPWR VPWR U$$2257/X sky130_fd_sc_hd__xor2_1
XU$$2268 U$$896/B1 U$$2308/A2 U$$3366/A1 U$$2308/B2 VGND VGND VPWR VPWR U$$2269/A
+ sky130_fd_sc_hd__a22o_1
XU$$1523 U$$1932/B1 U$$1557/A2 U$$1799/A1 U$$1557/B2 VGND VGND VPWR VPWR U$$1524/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2279 U$$2279/A U$$2317/B VGND VGND VPWR VPWR U$$2279/X sky130_fd_sc_hd__xor2_1
XU$$1534 U$$1534/A U$$1546/B VGND VGND VPWR VPWR U$$1534/X sky130_fd_sc_hd__xor2_1
XFILLER_163_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1545 U$$997/A1 U$$1545/A2 U$$997/B1 U$$1545/B2 VGND VGND VPWR VPWR U$$1546/A sky130_fd_sc_hd__a22o_1
XFILLER_76_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1556 U$$1556/A U$$1558/B VGND VGND VPWR VPWR U$$1556/X sky130_fd_sc_hd__xor2_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1567 U$$745/A1 U$$1591/A2 U$$610/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1568/A sky130_fd_sc_hd__a22o_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1578 U$$1578/A U$$1620/B VGND VGND VPWR VPWR U$$1578/X sky130_fd_sc_hd__xor2_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1589 U$$2683/B1 U$$1591/A2 U$$2550/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1590/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_108_0 dadda_fa_7_108_0/A dadda_fa_7_108_0/B dadda_fa_7_108_0/CIN VGND
+ VGND VPWR VPWR _405_/D _276_/D sky130_fd_sc_hd__fa_1
XFILLER_200_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_84_0_1854 VGND VGND VPWR VPWR dadda_fa_1_84_0/A dadda_fa_1_84_0_1854/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_111_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater401 U$$793/A2 VGND VGND VPWR VPWR U$$783/A2 sky130_fd_sc_hd__buf_4
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_1 dadda_fa_2_60_1/A dadda_fa_2_60_1/B dadda_fa_2_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_0/CIN dadda_fa_3_60_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_97_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$208 final_adder.U$$208/A final_adder.U$$208/B VGND VGND VPWR VPWR
+ final_adder.U$$336/B sky130_fd_sc_hd__and2_1
XFILLER_170_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater412 U$$678/A2 VGND VGND VPWR VPWR U$$636/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$219 final_adder.U$$218/B final_adder.U$$989/B1 final_adder.U$$219/B1
+ VGND VGND VPWR VPWR final_adder.U$$219/X sky130_fd_sc_hd__a21o_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater423 U$$527/A2 VGND VGND VPWR VPWR U$$473/A2 sky130_fd_sc_hd__buf_4
Xrepeater434 U$$4226/A2 VGND VGND VPWR VPWR U$$4210/A2 sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_2_53_0 dadda_fa_2_53_0/A dadda_fa_2_53_0/B dadda_fa_2_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_0/B dadda_fa_3_53_2/B sky130_fd_sc_hd__fa_1
XFILLER_211_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater445 U$$94/A2 VGND VGND VPWR VPWR U$$134/A2 sky130_fd_sc_hd__buf_8
XFILLER_84_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater456 U$$3874/A2 VGND VGND VPWR VPWR U$$3902/A2 sky130_fd_sc_hd__buf_6
XFILLER_66_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater467 U$$3777/A2 VGND VGND VPWR VPWR U$$3833/A2 sky130_fd_sc_hd__buf_6
Xrepeater478 U$$3566/X VGND VGND VPWR VPWR U$$3636/A2 sky130_fd_sc_hd__buf_4
XU$$4160 input78/X U$$4176/A2 U$$4162/A1 U$$4176/B2 VGND VGND VPWR VPWR U$$4161/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater489 U$$3378/A2 VGND VGND VPWR VPWR U$$3348/A2 sky130_fd_sc_hd__clkbuf_8
XU$$4171 U$$4171/A U$$4246/A VGND VGND VPWR VPWR U$$4171/X sky130_fd_sc_hd__xor2_1
XFILLER_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4182 U$$4456/A1 U$$4226/A2 input91/X U$$4226/B2 VGND VGND VPWR VPWR U$$4183/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_896 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4193 U$$4193/A U$$4211/B VGND VGND VPWR VPWR U$$4193/X sky130_fd_sc_hd__xor2_1
XFILLER_129_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3470 U$$3470/A U$$3504/B VGND VGND VPWR VPWR U$$3470/X sky130_fd_sc_hd__xor2_1
XFILLER_80_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3481 U$$3481/A1 U$$3489/A2 U$$741/B1 U$$3489/B2 VGND VGND VPWR VPWR U$$3482/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_1038 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3492 U$$3492/A U$$3518/B VGND VGND VPWR VPWR U$$3492/X sky130_fd_sc_hd__xor2_1
XFILLER_80_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_7_0 U$$21/X U$$154/X U$$287/X VGND VGND VPWR VPWR dadda_fa_6_8_0/A dadda_fa_6_7_0/CIN
+ sky130_fd_sc_hd__fa_1
XU$$2780 input72/X U$$2868/A2 U$$4013/B1 U$$2868/B2 VGND VGND VPWR VPWR U$$2781/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2791 U$$2791/A U$$2797/B VGND VGND VPWR VPWR U$$2791/X sky130_fd_sc_hd__xor2_1
XFILLER_90_1115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1787_1723 VGND VGND VPWR VPWR U$$1787_1723/HI U$$1787/A1 sky130_fd_sc_hd__conb_1
XFILLER_119_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_82_2 dadda_fa_4_82_2/A dadda_fa_4_82_2/B dadda_fa_4_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_83_0/CIN dadda_fa_5_82_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_75_1 dadda_fa_4_75_1/A dadda_fa_4_75_1/B dadda_fa_4_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/B dadda_fa_5_75_1/B sky130_fd_sc_hd__fa_1
XFILLER_150_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_52_0 dadda_fa_7_52_0/A dadda_fa_7_52_0/B dadda_fa_7_52_0/CIN VGND VGND
+ VPWR VPWR _349_/D _220_/D sky130_fd_sc_hd__fa_2
XFILLER_1_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_68_0 dadda_fa_4_68_0/A dadda_fa_4_68_0/B dadda_fa_4_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/A dadda_fa_5_68_1/A sky130_fd_sc_hd__fa_1
Xinput204 c[52] VGND VGND VPWR VPWR input204/X sky130_fd_sc_hd__buf_2
XFILLER_130_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput215 c[62] VGND VGND VPWR VPWR input215/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput226 c[72] VGND VGND VPWR VPWR input226/X sky130_fd_sc_hd__clkbuf_2
XTAP_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 c[82] VGND VGND VPWR VPWR input237/X sky130_fd_sc_hd__buf_2
XTAP_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput248 c[92] VGND VGND VPWR VPWR input248/X sky130_fd_sc_hd__clkbuf_4
XFILLER_88_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$720 final_adder.U$$720/A final_adder.U$$720/B VGND VGND VPWR VPWR
+ final_adder.U$$800/A sky130_fd_sc_hd__and2_1
XTAP_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$731 final_adder.U$$714/A final_adder.U$$503/X final_adder.U$$611/X
+ VGND VGND VPWR VPWR final_adder.U$$731/X sky130_fd_sc_hd__a21o_2
XTAP_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$742 final_adder.U$$774/B final_adder.U$$742/B VGND VGND VPWR VPWR
+ final_adder.U$$742/X sky130_fd_sc_hd__and2_1
XTAP_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$753 final_adder.U$$752/B final_adder.U$$673/X final_adder.U$$641/X
+ VGND VGND VPWR VPWR final_adder.U$$753/X sky130_fd_sc_hd__a21o_1
XTAP_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$764 final_adder.U$$796/B final_adder.U$$764/B VGND VGND VPWR VPWR
+ final_adder.U$$764/X sky130_fd_sc_hd__and2_1
XFILLER_5_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$603 U$$603/A U$$637/B VGND VGND VPWR VPWR U$$603/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$775 final_adder.U$$774/B final_adder.U$$695/X final_adder.U$$663/X
+ VGND VGND VPWR VPWR final_adder.U$$775/X sky130_fd_sc_hd__a21o_1
XU$$614 U$$66/A1 U$$616/A2 U$$68/A1 U$$616/B2 VGND VGND VPWR VPWR U$$615/A sky130_fd_sc_hd__a22o_1
XFILLER_72_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$786 final_adder.U$$786/A final_adder.U$$786/B VGND VGND VPWR VPWR
+ final_adder.U$$786/X sky130_fd_sc_hd__and2_1
XFILLER_29_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater990 U$$1209/B VGND VGND VPWR VPWR U$$1205/B sky130_fd_sc_hd__buf_6
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$625 U$$625/A U$$625/B VGND VGND VPWR VPWR U$$625/X sky130_fd_sc_hd__xor2_1
XFILLER_72_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$797 final_adder.U$$796/B final_adder.U$$717/X final_adder.U$$685/X
+ VGND VGND VPWR VPWR final_adder.U$$797/X sky130_fd_sc_hd__a21o_1
XFILLER_72_833 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$636 U$$910/A1 U$$636/A2 U$$773/B1 U$$636/B2 VGND VGND VPWR VPWR U$$637/A sky130_fd_sc_hd__a22o_1
XFILLER_205_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$647 U$$647/A U$$651/B VGND VGND VPWR VPWR U$$647/X sky130_fd_sc_hd__xor2_1
XFILLER_147_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$658 U$$930/B1 U$$678/A2 U$$660/A1 U$$678/B2 VGND VGND VPWR VPWR U$$659/A sky130_fd_sc_hd__a22o_1
XFILLER_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$669 U$$669/A U$$673/B VGND VGND VPWR VPWR U$$669/X sky130_fd_sc_hd__xor2_1
XFILLER_72_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_500 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1503 U$$3555/B1 VGND VGND VPWR VPWR U$$4103/B1 sky130_fd_sc_hd__buf_4
Xrepeater1514 U$$950/A1 VGND VGND VPWR VPWR U$$2044/B1 sky130_fd_sc_hd__buf_6
Xrepeater1525 U$$3852/B1 VGND VGND VPWR VPWR U$$2621/A1 sky130_fd_sc_hd__buf_4
Xrepeater1536 U$$3/A VGND VGND VPWR VPWR U$$99/B sky130_fd_sc_hd__buf_8
XFILLER_4_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1547 U$$946/A1 VGND VGND VPWR VPWR U$$944/B1 sky130_fd_sc_hd__buf_6
Xrepeater1558 U$$2312/B1 VGND VGND VPWR VPWR U$$807/A1 sky130_fd_sc_hd__buf_4
Xrepeater1569 U$$4504/A1 VGND VGND VPWR VPWR U$$4365/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_3_70_0 dadda_fa_3_70_0/A dadda_fa_3_70_0/B dadda_fa_3_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_0/B dadda_fa_4_70_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2010 U$$2967/B1 U$$2046/A2 U$$2834/A1 U$$2046/B2 VGND VGND VPWR VPWR U$$2011/A
+ sky130_fd_sc_hd__a22o_1
XU$$2021 U$$2021/A U$$2054/A VGND VGND VPWR VPWR U$$2021/X sky130_fd_sc_hd__xor2_1
XFILLER_62_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2032 U$$2032/A1 U$$2046/A2 U$$936/B1 U$$2046/B2 VGND VGND VPWR VPWR U$$2033/A
+ sky130_fd_sc_hd__a22o_1
XU$$2043 U$$2043/A U$$2043/B VGND VGND VPWR VPWR U$$2043/X sky130_fd_sc_hd__xor2_1
XU$$2054 U$$2054/A VGND VGND VPWR VPWR U$$2054/Y sky130_fd_sc_hd__inv_1
XU$$2065 U$$2202/A1 U$$2093/A2 U$$2065/B1 U$$2093/B2 VGND VGND VPWR VPWR U$$2066/A
+ sky130_fd_sc_hd__a22o_1
XU$$1320 U$$1320/A U$$1354/B VGND VGND VPWR VPWR U$$1320/X sky130_fd_sc_hd__xor2_1
XU$$1331 U$$2975/A1 U$$1337/A2 U$$2975/B1 U$$1337/B2 VGND VGND VPWR VPWR U$$1332/A
+ sky130_fd_sc_hd__a22o_1
XU$$2076 U$$2076/A U$$2094/B VGND VGND VPWR VPWR U$$2076/X sky130_fd_sc_hd__xor2_1
XFILLER_204_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2087 U$$3594/A1 U$$2091/A2 U$$4005/B1 U$$2091/B2 VGND VGND VPWR VPWR U$$2088/A
+ sky130_fd_sc_hd__a22o_1
XU$$1342 U$$1342/A U$$1370/A VGND VGND VPWR VPWR U$$1342/X sky130_fd_sc_hd__xor2_1
XU$$2098 U$$2098/A U$$2100/B VGND VGND VPWR VPWR U$$2098/X sky130_fd_sc_hd__xor2_1
XU$$1353 U$$942/A1 U$$1353/A2 U$$944/A1 U$$1355/B2 VGND VGND VPWR VPWR U$$1354/A sky130_fd_sc_hd__a22o_1
XU$$1364 U$$1364/A U$$1366/B VGND VGND VPWR VPWR U$$1364/X sky130_fd_sc_hd__xor2_1
XFILLER_95_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1375 U$$1373/B input11/X input13/X U$$1370/Y VGND VGND VPWR VPWR U$$1375/X sky130_fd_sc_hd__a22o_4
XU$$1386 U$$1932/B1 U$$1422/A2 U$$1799/A1 U$$1422/B2 VGND VGND VPWR VPWR U$$1387/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1397 U$$1397/A U$$1399/B VGND VGND VPWR VPWR U$$1397/X sky130_fd_sc_hd__xor2_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_92_1 dadda_fa_5_92_1/A dadda_fa_5_92_1/B dadda_fa_5_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_93_0/B dadda_fa_7_92_0/A sky130_fd_sc_hd__fa_1
XFILLER_159_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_85_0 dadda_fa_5_85_0/A dadda_fa_5_85_0/B dadda_fa_5_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_86_0/A dadda_fa_6_85_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_190_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_77_7 U$$4151/X U$$4284/X U$$4417/X VGND VGND VPWR VPWR dadda_fa_2_78_2/CIN
+ dadda_fa_2_77_5/CIN sky130_fd_sc_hd__fa_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$60 _356_/Q _228_/Q VGND VGND VPWR VPWR final_adder.U$$965/B1 final_adder.U$$194/A
+ sky130_fd_sc_hd__ha_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$71 _367_/Q _239_/Q VGND VGND VPWR VPWR final_adder.U$$185/B1 final_adder.U$$184/B
+ sky130_fd_sc_hd__ha_1
XFILLER_54_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$82 _378_/Q _250_/Q VGND VGND VPWR VPWR final_adder.U$$943/B1 final_adder.U$$172/A
+ sky130_fd_sc_hd__ha_1
XFILLER_81_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$93 _389_/Q _261_/Q VGND VGND VPWR VPWR final_adder.U$$163/B1 final_adder.U$$162/B
+ sky130_fd_sc_hd__ha_1
XFILLER_81_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_101_2 dadda_fa_3_101_2/A dadda_fa_3_101_2/B dadda_fa_3_101_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_102_1/A dadda_fa_4_101_2/B sky130_fd_sc_hd__fa_1
XFILLER_107_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2737_1737 VGND VGND VPWR VPWR U$$2737_1737/HI U$$2737/B1 sky130_fd_sc_hd__conb_1
XFILLER_122_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_65_5 U$$2132/X U$$2265/X U$$2398/X VGND VGND VPWR VPWR dadda_fa_1_66_7/A
+ dadda_fa_2_65_0/A sky130_fd_sc_hd__fa_2
XTAP_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_115_0 dadda_fa_6_115_0/A dadda_fa_6_115_0/B dadda_fa_6_115_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_116_0/B dadda_fa_7_115_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$550 final_adder.U$$558/B final_adder.U$$550/B VGND VGND VPWR VPWR
+ final_adder.U$$670/B sky130_fd_sc_hd__and2_1
XTAP_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$561 final_adder.U$$560/B final_adder.U$$445/X final_adder.U$$437/X
+ VGND VGND VPWR VPWR final_adder.U$$561/X sky130_fd_sc_hd__a21o_1
XTAP_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$400 U$$674/A1 U$$278/X U$$676/A1 U$$279/X VGND VGND VPWR VPWR U$$401/A sky130_fd_sc_hd__a22o_1
XFILLER_45_811 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$572 final_adder.U$$580/B final_adder.U$$572/B VGND VGND VPWR VPWR
+ final_adder.U$$692/B sky130_fd_sc_hd__and2_1
XTAP_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$411 U$$411/A VGND VGND VPWR VPWR U$$411/Y sky130_fd_sc_hd__inv_1
XFILLER_205_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$583 final_adder.U$$582/B final_adder.U$$467/X final_adder.U$$459/X
+ VGND VGND VPWR VPWR final_adder.U$$583/X sky130_fd_sc_hd__a21o_1
XTAP_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$422 U$$422/A U$$436/B VGND VGND VPWR VPWR U$$422/X sky130_fd_sc_hd__xor2_1
XTAP_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_35_3 dadda_fa_3_35_3/A dadda_fa_3_35_3/B dadda_fa_3_35_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_36_1/B dadda_fa_4_35_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$594 final_adder.U$$602/B final_adder.U$$594/B VGND VGND VPWR VPWR
+ final_adder.U$$714/B sky130_fd_sc_hd__and2_1
XU$$433 U$$842/B1 U$$437/A2 U$$24/A1 U$$437/B2 VGND VGND VPWR VPWR U$$434/A sky130_fd_sc_hd__a22o_1
XTAP_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$444 U$$444/A U$$516/B VGND VGND VPWR VPWR U$$444/X sky130_fd_sc_hd__xor2_1
XFILLER_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$455 U$$864/B1 U$$491/A2 U$$731/A1 U$$491/B2 VGND VGND VPWR VPWR U$$456/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_28_2 dadda_fa_3_28_2/A dadda_fa_3_28_2/B dadda_fa_3_28_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_29_1/A dadda_fa_4_28_2/B sky130_fd_sc_hd__fa_1
XTAP_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$466 U$$466/A U$$484/B VGND VGND VPWR VPWR U$$466/X sky130_fd_sc_hd__xor2_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$477 U$$477/A1 U$$527/A2 U$$68/A1 U$$527/B2 VGND VGND VPWR VPWR U$$478/A sky130_fd_sc_hd__a22o_1
XFILLER_205_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$488 U$$488/A U$$492/B VGND VGND VPWR VPWR U$$488/X sky130_fd_sc_hd__xor2_1
XU$$499 U$$910/A1 U$$527/A2 U$$773/B1 U$$527/B2 VGND VGND VPWR VPWR U$$500/A sky130_fd_sc_hd__a22o_1
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_587 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_982 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1300 U$$3510/B VGND VGND VPWR VPWR U$$3504/B sky130_fd_sc_hd__buf_6
Xrepeater1311 input44/X VGND VGND VPWR VPWR U$$3377/B sky130_fd_sc_hd__buf_6
XFILLER_158_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1322 U$$3077/B VGND VGND VPWR VPWR U$$3075/B sky130_fd_sc_hd__buf_8
XFILLER_201_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1333 U$$2968/B VGND VGND VPWR VPWR U$$2950/B sky130_fd_sc_hd__buf_6
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1344 U$$2859/B VGND VGND VPWR VPWR U$$2869/B sky130_fd_sc_hd__buf_6
Xrepeater1355 U$$272/B VGND VGND VPWR VPWR U$$260/B sky130_fd_sc_hd__buf_6
XFILLER_125_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1366 U$$2601/B VGND VGND VPWR VPWR U$$2597/B sky130_fd_sc_hd__buf_6
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1377 U$$794/B VGND VGND VPWR VPWR U$$770/B sky130_fd_sc_hd__buf_8
Xrepeater1388 U$$2466/A VGND VGND VPWR VPWR U$$2446/B sky130_fd_sc_hd__buf_8
XFILLER_113_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1399 input27/X VGND VGND VPWR VPWR U$$2303/B sky130_fd_sc_hd__buf_6
XFILLER_84_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_1264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_2_31_4 U$$1665/X U$$1798/X VGND VGND VPWR VPWR dadda_fa_3_32_2/A dadda_fa_4_31_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_122_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_7_1_0 U$$9/X input168/X VGND VGND VPWR VPWR _298_/D _169_/D sky130_fd_sc_hd__ha_1
XFILLER_48_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_30_2 U$$865/X U$$998/X U$$1131/X VGND VGND VPWR VPWR dadda_fa_3_31_1/CIN
+ dadda_fa_3_30_3/B sky130_fd_sc_hd__fa_1
XFILLER_211_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1150 U$$328/A1 U$$1162/A2 U$$328/B1 U$$1162/B2 VGND VGND VPWR VPWR U$$1151/A sky130_fd_sc_hd__a22o_1
XFILLER_211_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1161 U$$1161/A U$$1205/B VGND VGND VPWR VPWR U$$1161/X sky130_fd_sc_hd__xor2_1
XU$$1172 U$$1446/A1 U$$1174/A2 U$$1448/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1173/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1183 U$$1183/A U$$1223/B VGND VGND VPWR VPWR U$$1183/X sky130_fd_sc_hd__xor2_1
XU$$1194 U$$98/A1 U$$1204/A2 U$$98/B1 U$$1204/B2 VGND VGND VPWR VPWR U$$1195/A sky130_fd_sc_hd__a22o_1
XFILLER_148_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_82_5 U$$3230/X U$$3363/X U$$3496/X VGND VGND VPWR VPWR dadda_fa_2_83_3/A
+ dadda_fa_2_82_5/B sky130_fd_sc_hd__fa_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_75_4 U$$3216/X U$$3349/X U$$3482/X VGND VGND VPWR VPWR dadda_fa_2_76_1/CIN
+ dadda_fa_2_75_4/CIN sky130_fd_sc_hd__fa_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_3 U$$3734/X U$$3867/X U$$4000/X VGND VGND VPWR VPWR dadda_fa_2_69_1/B
+ dadda_fa_2_68_4/B sky130_fd_sc_hd__fa_1
XFILLER_112_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_45_2 dadda_fa_4_45_2/A dadda_fa_4_45_2/B dadda_fa_4_45_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_46_0/CIN dadda_fa_5_45_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_1 dadda_fa_4_38_1/A dadda_fa_4_38_1/B dadda_fa_4_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/B dadda_fa_5_38_1/B sky130_fd_sc_hd__fa_1
XFILLER_100_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_15_0 dadda_fa_7_15_0/A dadda_fa_7_15_0/B dadda_fa_7_15_0/CIN VGND VGND
+ VPWR VPWR _312_/D _183_/D sky130_fd_sc_hd__fa_1
XFILLER_148_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_106 _384_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_117 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_128 _420_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 U$$3082/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ _411_/CLK _280_/D VGND VGND VPWR VPWR _280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_418 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2600_1734 VGND VGND VPWR VPWR U$$2600_1734/HI U$$2600/B1 sky130_fd_sc_hd__conb_1
XFILLER_5_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_700 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_70_3 U$$1610/X U$$1743/X U$$1876/X VGND VGND VPWR VPWR dadda_fa_1_71_7/B
+ dadda_fa_1_70_8/CIN sky130_fd_sc_hd__fa_1
XTAP_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_2 U$$931/X U$$1064/X U$$1197/X VGND VGND VPWR VPWR dadda_fa_1_64_6/A
+ dadda_fa_1_63_8/A sky130_fd_sc_hd__fa_1
XFILLER_77_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_40_1 dadda_fa_3_40_1/A dadda_fa_3_40_1/B dadda_fa_3_40_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_0/CIN dadda_fa_4_40_2/A sky130_fd_sc_hd__fa_1
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_56_1 U$$518/X U$$651/X U$$784/X VGND VGND VPWR VPWR dadda_fa_1_57_7/CIN
+ dadda_fa_1_56_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_56_clk clkbuf_3_1_0_clk/X VGND VGND VPWR VPWR _363_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_33_0 input183/X dadda_fa_3_33_0/B dadda_fa_3_33_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_34_0/B dadda_fa_4_33_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$230 U$$230/A U$$264/B VGND VGND VPWR VPWR U$$230/X sky130_fd_sc_hd__xor2_1
XFILLER_45_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$391 final_adder.U$$390/B final_adder.U$$269/X final_adder.U$$265/X
+ VGND VGND VPWR VPWR final_adder.U$$391/X sky130_fd_sc_hd__a21o_2
XTAP_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$241 U$$926/A1 U$$243/A2 U$$654/A1 U$$243/B2 VGND VGND VPWR VPWR U$$242/A sky130_fd_sc_hd__a22o_1
XTAP_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$252 U$$252/A U$$260/B VGND VGND VPWR VPWR U$$252/X sky130_fd_sc_hd__xor2_1
XFILLER_206_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$263 U$$674/A1 U$$263/A2 U$$676/A1 U$$142/X VGND VGND VPWR VPWR U$$264/A sky130_fd_sc_hd__a22o_1
XFILLER_72_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$274 U$$274/A VGND VGND VPWR VPWR U$$274/Y sky130_fd_sc_hd__inv_1
XFILLER_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$285 U$$285/A U$$317/B VGND VGND VPWR VPWR U$$285/X sky130_fd_sc_hd__xor2_1
XU$$296 U$$842/B1 U$$302/A2 U$$24/A1 U$$302/B2 VGND VGND VPWR VPWR U$$297/A sky130_fd_sc_hd__a22o_1
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2 U$$3/A VGND VGND VPWR VPWR U$$2/Y sky130_fd_sc_hd__inv_1
XFILLER_69_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput305 output305/A VGND VGND VPWR VPWR o[28] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_4 input248/X dadda_fa_2_92_4/B dadda_fa_2_92_4/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_93_1/CIN dadda_fa_3_92_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1130 U$$40/A1 VGND VGND VPWR VPWR U$$999/A1 sky130_fd_sc_hd__buf_6
XFILLER_58_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput316 output316/A VGND VGND VPWR VPWR o[38] sky130_fd_sc_hd__buf_2
Xoutput327 output327/A VGND VGND VPWR VPWR o[48] sky130_fd_sc_hd__buf_2
XFILLER_142_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1141 U$$4011/A1 VGND VGND VPWR VPWR U$$721/B1 sky130_fd_sc_hd__buf_6
Xoutput338 output338/A VGND VGND VPWR VPWR o[58] sky130_fd_sc_hd__buf_2
Xrepeater1152 U$$4146/A1 VGND VGND VPWR VPWR U$$4144/B1 sky130_fd_sc_hd__buf_12
Xoutput349 output349/A VGND VGND VPWR VPWR o[68] sky130_fd_sc_hd__buf_2
Xrepeater1163 U$$32/B1 VGND VGND VPWR VPWR U$$34/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_85_3 dadda_fa_2_85_3/A dadda_fa_2_85_3/B dadda_fa_2_85_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/B dadda_fa_3_85_3/B sky130_fd_sc_hd__fa_1
XFILLER_153_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1174 U$$4005/A1 VGND VGND VPWR VPWR U$$3594/A1 sky130_fd_sc_hd__buf_4
Xrepeater1185 U$$3727/B1 VGND VGND VPWR VPWR U$$2357/B1 sky130_fd_sc_hd__buf_4
XFILLER_102_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1196 input66/X VGND VGND VPWR VPWR U$$4410/B1 sky130_fd_sc_hd__buf_8
XFILLER_113_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_78_2 dadda_fa_2_78_2/A dadda_fa_2_78_2/B dadda_fa_2_78_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/A dadda_fa_3_78_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_55_1 dadda_fa_5_55_1/A dadda_fa_5_55_1/B dadda_fa_5_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_56_0/B dadda_fa_7_55_0/A sky130_fd_sc_hd__fa_1
XFILLER_68_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_48_0 dadda_fa_5_48_0/A dadda_fa_5_48_0/B dadda_fa_5_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_49_0/A dadda_fa_6_48_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_2_22_0 U$$51/X U$$184/X VGND VGND VPWR VPWR dadda_fa_3_23_3/CIN dadda_fa_4_22_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_55_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_101_1 U$$3002/X U$$3135/X U$$3268/X VGND VGND VPWR VPWR dadda_fa_3_102_2/A
+ dadda_fa_3_101_3/B sky130_fd_sc_hd__fa_1
XFILLER_36_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_122_0 U$$4241/X U$$4374/X U$$4507/X VGND VGND VPWR VPWR dadda_fa_6_123_0/A
+ dadda_fa_6_122_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_80_2 U$$1896/X U$$2029/X U$$2162/X VGND VGND VPWR VPWR dadda_fa_2_81_1/B
+ dadda_fa_2_80_4/A sky130_fd_sc_hd__fa_1
XFILLER_104_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_73_1 U$$2281/X U$$2414/X U$$2547/X VGND VGND VPWR VPWR dadda_fa_2_74_0/CIN
+ dadda_fa_2_73_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_50_0 dadda_fa_4_50_0/A dadda_fa_4_50_0/B dadda_fa_4_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/A dadda_fa_5_50_1/A sky130_fd_sc_hd__fa_1
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_66_0 U$$2533/X U$$2666/X U$$2799/X VGND VGND VPWR VPWR dadda_fa_2_67_0/B
+ dadda_fa_2_66_3/B sky130_fd_sc_hd__fa_1
XFILLER_150_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4413_1783 VGND VGND VPWR VPWR U$$4413_1783/HI U$$4413/B sky130_fd_sc_hd__conb_1
XFILLER_86_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2609 U$$2609/A1 U$$2625/A2 U$$2609/B1 U$$2625/B2 VGND VGND VPWR VPWR U$$2610/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk _239_/CLK VGND VGND VPWR VPWR _376_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1908 U$$1908/A U$$1912/B VGND VGND VPWR VPWR U$$1908/X sky130_fd_sc_hd__xor2_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_401_ _401_/CLK _401_/D VGND VGND VPWR VPWR _401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1919 input21/X VGND VGND VPWR VPWR U$$1921/B sky130_fd_sc_hd__inv_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_332_ _342_/CLK _332_/D VGND VGND VPWR VPWR _332_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_830 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_263_ _390_/CLK _263_/D VGND VGND VPWR VPWR _263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_194_ _323_/CLK _194_/D VGND VGND VPWR VPWR _194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_95_2 dadda_fa_3_95_2/A dadda_fa_3_95_2/B dadda_fa_3_95_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_1/A dadda_fa_4_95_2/B sky130_fd_sc_hd__fa_1
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_88_1 dadda_fa_3_88_1/A dadda_fa_3_88_1/B dadda_fa_3_88_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_0/CIN dadda_fa_4_88_2/A sky130_fd_sc_hd__fa_1
XFILLER_123_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_65_0 dadda_fa_6_65_0/A dadda_fa_6_65_0/B dadda_fa_6_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_66_0/B dadda_fa_7_65_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1045 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater808 U$$2302/B2 VGND VGND VPWR VPWR U$$2252/B2 sky130_fd_sc_hd__clkbuf_8
Xrepeater819 U$$2183/B2 VGND VGND VPWR VPWR U$$2189/B2 sky130_fd_sc_hd__buf_6
XU$$4501 U$$4501/A U$$4501/B VGND VGND VPWR VPWR U$$4501/X sky130_fd_sc_hd__xor2_1
XU$$4512 U$$4512/A1 U$$4388/X U$$4514/A1 U$$4512/B2 VGND VGND VPWR VPWR U$$4513/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3800 U$$3800/A U$$3814/B VGND VGND VPWR VPWR U$$3800/X sky130_fd_sc_hd__xor2_1
XU$$15 U$$15/A U$$9/B VGND VGND VPWR VPWR U$$15/X sky130_fd_sc_hd__xor2_1
XU$$3811 U$$3946/B1 U$$3813/A2 U$$3813/A1 U$$3813/B2 VGND VGND VPWR VPWR U$$3812/A
+ sky130_fd_sc_hd__a22o_1
XU$$26 U$$26/A1 U$$8/A2 U$$28/A1 U$$8/B2 VGND VGND VPWR VPWR U$$27/A sky130_fd_sc_hd__a22o_1
XTAP_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_747 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3822 U$$3822/A U$$3826/B VGND VGND VPWR VPWR U$$3822/X sky130_fd_sc_hd__xor2_1
XU$$37 U$$37/A U$$43/B VGND VGND VPWR VPWR U$$37/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_117_1 U$$4098/X U$$4231/X U$$4364/X VGND VGND VPWR VPWR dadda_fa_5_118_0/B
+ dadda_fa_5_117_1/B sky130_fd_sc_hd__fa_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_clk _255_/CLK VGND VGND VPWR VPWR _420_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3833 U$$4242/B1 U$$3833/A2 U$$3833/B1 U$$3833/B2 VGND VGND VPWR VPWR U$$3834/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$48 U$$48/A1 U$$50/A2 U$$48/B1 U$$50/B2 VGND VGND VPWR VPWR U$$49/A sky130_fd_sc_hd__a22o_1
XU$$3844 U$$3979/B1 U$$3878/A2 U$$832/A1 U$$3878/B2 VGND VGND VPWR VPWR U$$3845/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$59 U$$59/A U$$85/B VGND VGND VPWR VPWR U$$59/X sky130_fd_sc_hd__xor2_1
XU$$3855 U$$3855/A U$$3875/B VGND VGND VPWR VPWR U$$3855/X sky130_fd_sc_hd__xor2_1
XTAP_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3866 U$$4275/B1 U$$3902/A2 U$$4277/B1 U$$3902/B2 VGND VGND VPWR VPWR U$$3867/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3877 U$$3877/A U$$3879/B VGND VGND VPWR VPWR U$$3877/X sky130_fd_sc_hd__xor2_1
XTAP_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3888 input79/X U$$3970/A2 input80/X U$$3970/B2 VGND VGND VPWR VPWR U$$3889/A sky130_fd_sc_hd__a22o_1
XTAP_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3899 U$$3899/A U$$3903/B VGND VGND VPWR VPWR U$$3899/X sky130_fd_sc_hd__xor2_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_17 _329_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _337_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_39 _340_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_90_1 U$$3645/X U$$3778/X U$$3911/X VGND VGND VPWR VPWR dadda_fa_3_91_0/CIN
+ dadda_fa_3_90_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_115_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_83_0 U$$4163/X U$$4296/X U$$4429/X VGND VGND VPWR VPWR dadda_fa_3_84_0/B
+ dadda_fa_3_83_2/B sky130_fd_sc_hd__fa_1
XFILLER_142_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_52_6 U$$2771/X U$$2904/X U$$3037/X VGND VGND VPWR VPWR dadda_fa_2_53_2/B
+ dadda_fa_2_52_5/B sky130_fd_sc_hd__fa_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_4_0 dadda_fa_7_4_0/A dadda_fa_7_4_0/B dadda_fa_7_4_0/CIN VGND VGND VPWR
+ VPWR _301_/D _172_/D sky130_fd_sc_hd__fa_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4443_1798 VGND VGND VPWR VPWR U$$4443_1798/HI U$$4443/B sky130_fd_sc_hd__conb_1
XFILLER_211_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1009 final_adder.U$$238/A final_adder.U$$619/X final_adder.U$$239/A2
+ VGND VGND VPWR VPWR final_adder.U$$1041/B sky130_fd_sc_hd__a21o_1
XFILLER_164_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_82_0 dadda_fa_7_82_0/A dadda_fa_7_82_0/B dadda_fa_7_82_0/CIN VGND VGND
+ VPWR VPWR _379_/D _250_/D sky130_fd_sc_hd__fa_2
Xdadda_fa_4_98_0 dadda_fa_4_98_0/A dadda_fa_4_98_0/B dadda_fa_4_98_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/A dadda_fa_5_98_1/A sky130_fd_sc_hd__fa_1
XFILLER_194_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1067 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_76 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1040 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3107 U$$3107/A U$$3109/B VGND VGND VPWR VPWR U$$3107/X sky130_fd_sc_hd__xor2_1
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3118 U$$789/A1 U$$3118/A2 U$$517/A1 U$$3118/B2 VGND VGND VPWR VPWR U$$3119/A sky130_fd_sc_hd__a22o_1
XFILLER_46_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3129 U$$3129/A U$$3133/B VGND VGND VPWR VPWR U$$3129/X sky130_fd_sc_hd__xor2_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2406 U$$2406/A U$$2446/B VGND VGND VPWR VPWR U$$2406/X sky130_fd_sc_hd__xor2_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1504_1718 VGND VGND VPWR VPWR U$$1504_1718/HI U$$1504/B1 sky130_fd_sc_hd__conb_1
XFILLER_62_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2417 U$$3922/B1 U$$2417/A2 U$$3787/B1 U$$2417/B2 VGND VGND VPWR VPWR U$$2418/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2428 U$$2428/A U$$2454/B VGND VGND VPWR VPWR U$$2428/X sky130_fd_sc_hd__xor2_1
XU$$2439 U$$2711/B1 U$$2333/X U$$934/A1 U$$2334/X VGND VGND VPWR VPWR U$$2440/A sky130_fd_sc_hd__a22o_1
XFILLER_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1705 U$$1705/A U$$1707/B VGND VGND VPWR VPWR U$$1705/X sky130_fd_sc_hd__xor2_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1716 U$$4456/A1 U$$1764/A2 U$$2951/A1 U$$1764/B2 VGND VGND VPWR VPWR U$$1717/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_633 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1727 U$$1727/A U$$1739/B VGND VGND VPWR VPWR U$$1727/X sky130_fd_sc_hd__xor2_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1738 U$$3108/A1 U$$1746/A2 U$$2425/A1 U$$1746/B2 VGND VGND VPWR VPWR U$$1739/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1749 U$$1749/A U$$1765/B VGND VGND VPWR VPWR U$$1749/X sky130_fd_sc_hd__xor2_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_315_ _326_/CLK _315_/D VGND VGND VPWR VPWR _315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_246_ _246_/CLK _246_/D VGND VGND VPWR VPWR _246_/Q sky130_fd_sc_hd__dfxtp_1
Xinput15 a[22] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput26 a[32] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput37 a[42] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 a[52] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput59 a[62] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_1
X_177_ _326_/CLK _177_/D VGND VGND VPWR VPWR _177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_62_5 dadda_fa_2_62_5/A dadda_fa_2_62_5/B dadda_fa_2_62_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_63_2/A dadda_fa_4_62_0/A sky130_fd_sc_hd__fa_2
XFILLER_111_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater605 U$$1607/A2 VGND VGND VPWR VPWR U$$1591/A2 sky130_fd_sc_hd__buf_6
XFILLER_111_468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater616 U$$1502/A2 VGND VGND VPWR VPWR U$$1448/A2 sky130_fd_sc_hd__buf_4
Xrepeater627 U$$1289/A2 VGND VGND VPWR VPWR U$$1271/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_55_4 dadda_fa_2_55_4/A dadda_fa_2_55_4/B dadda_fa_2_55_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_1/CIN dadda_fa_3_55_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater638 U$$1204/A2 VGND VGND VPWR VPWR U$$1162/A2 sky130_fd_sc_hd__buf_4
XU$$4320 U$$4320/A U$$4330/B VGND VGND VPWR VPWR U$$4320/X sky130_fd_sc_hd__xor2_1
Xrepeater649 U$$892/B2 VGND VGND VPWR VPWR U$$882/B2 sky130_fd_sc_hd__buf_4
XU$$4331 U$$4466/B1 U$$4349/A2 U$$4333/A1 U$$4349/B2 VGND VGND VPWR VPWR U$$4332/A
+ sky130_fd_sc_hd__a22o_1
XU$$4342 U$$4342/A U$$4354/B VGND VGND VPWR VPWR U$$4342/X sky130_fd_sc_hd__xor2_1
XFILLER_77_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4353 U$$4490/A1 U$$4361/A2 U$$4492/A1 U$$4361/B2 VGND VGND VPWR VPWR U$$4354/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4364 U$$4364/A input60/X VGND VGND VPWR VPWR U$$4364/X sky130_fd_sc_hd__xor2_1
XFILLER_38_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_48_3 dadda_fa_2_48_3/A dadda_fa_2_48_3/B dadda_fa_2_48_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/B dadda_fa_3_48_3/B sky130_fd_sc_hd__fa_1
XU$$3630 U$$4176/B1 U$$3636/A2 U$$4043/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3631/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4375 U$$4512/A1 U$$4251/X U$$4375/B1 U$$4252/X VGND VGND VPWR VPWR U$$4376/A sky130_fd_sc_hd__a22o_1
XU$$4386 U$$4386/A VGND VGND VPWR VPWR U$$4386/Y sky130_fd_sc_hd__inv_1
XU$$3641 U$$3641/A U$$3643/B VGND VGND VPWR VPWR U$$3641/X sky130_fd_sc_hd__xor2_1
XU$$3652 U$$3787/B1 U$$3680/A2 U$$4476/A1 U$$3680/B2 VGND VGND VPWR VPWR U$$3653/A
+ sky130_fd_sc_hd__a22o_1
XU$$4397 U$$4397/A U$$4397/B VGND VGND VPWR VPWR U$$4397/X sky130_fd_sc_hd__xor2_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3663 U$$3663/A U$$3665/B VGND VGND VPWR VPWR U$$3663/X sky130_fd_sc_hd__xor2_1
XU$$3674 U$$3946/B1 U$$3680/A2 U$$3813/A1 U$$3680/B2 VGND VGND VPWR VPWR U$$3675/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2940 U$$2940/A U$$2968/B VGND VGND VPWR VPWR U$$2940/X sky130_fd_sc_hd__xor2_1
XU$$3685 U$$3685/A U$$3698/A VGND VGND VPWR VPWR U$$3685/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_18_1 dadda_fa_5_18_1/A dadda_fa_5_18_1/B dadda_fa_5_18_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_19_0/B dadda_fa_7_18_0/A sky130_fd_sc_hd__fa_1
XU$$2951 U$$2951/A1 U$$2995/A2 U$$2951/B1 U$$2995/B2 VGND VGND VPWR VPWR U$$2952/A
+ sky130_fd_sc_hd__a22o_1
XU$$3696 U$$4242/B1 U$$3696/A2 U$$3696/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3697/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2962 U$$2962/A U$$3008/B VGND VGND VPWR VPWR U$$2962/X sky130_fd_sc_hd__xor2_1
XU$$2973 U$$3108/B1 U$$2977/A2 U$$2975/A1 U$$2979/B2 VGND VGND VPWR VPWR U$$2974/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2984 U$$2984/A U$$3008/B VGND VGND VPWR VPWR U$$2984/X sky130_fd_sc_hd__xor2_1
XU$$2995 U$$392/A1 U$$2995/A2 U$$3545/A1 U$$2995/B2 VGND VGND VPWR VPWR U$$2996/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_636 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_9_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _337_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$913 final_adder.U$$142/A final_adder.U$$851/X final_adder.U$$913/B1
+ VGND VGND VPWR VPWR final_adder.U$$913/X sky130_fd_sc_hd__a21o_1
XTAP_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$935 final_adder.U$$164/A ANTENNA_250/DIODE final_adder.U$$935/B1 VGND
+ VGND VPWR VPWR final_adder.U$$935/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_3 U$$1304/X U$$1437/X U$$1570/X VGND VGND VPWR VPWR dadda_fa_2_51_1/B
+ dadda_fa_2_50_4/B sky130_fd_sc_hd__fa_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$957 final_adder.U$$186/A final_adder.U$$895/X final_adder.U$$957/B1
+ VGND VGND VPWR VPWR final_adder.U$$957/X sky130_fd_sc_hd__a21o_1
XU$$807 U$$807/A1 U$$689/X U$$807/B1 U$$690/X VGND VGND VPWR VPWR U$$808/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$979 final_adder.U$$208/A final_adder.U$$821/X final_adder.U$$979/B1
+ VGND VGND VPWR VPWR final_adder.U$$979/X sky130_fd_sc_hd__a21o_1
XU$$818 U$$818/A U$$821/A VGND VGND VPWR VPWR U$$818/X sky130_fd_sc_hd__xor2_1
XU$$829 U$$829/A U$$919/B VGND VGND VPWR VPWR U$$829/X sky130_fd_sc_hd__xor2_1
XFILLER_16_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_43_2 U$$891/X U$$1024/X U$$1157/X VGND VGND VPWR VPWR dadda_fa_2_44_3/B
+ dadda_fa_2_43_5/B sky130_fd_sc_hd__fa_1
XFILLER_95_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_20_1 dadda_fa_4_20_1/A dadda_fa_4_20_1/B dadda_fa_4_20_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_21_0/B dadda_fa_5_20_1/B sky130_fd_sc_hd__fa_1
XFILLER_37_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3833_1754 VGND VGND VPWR VPWR U$$3833_1754/HI U$$3833/B1 sky130_fd_sc_hd__conb_1
XFILLER_197_700 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_13_0 U$$33/X U$$166/X U$$299/X VGND VGND VPWR VPWR dadda_fa_5_14_0/A dadda_fa_5_13_1/A
+ sky130_fd_sc_hd__fa_1
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1707 U$$4335/B1 VGND VGND VPWR VPWR U$$3787/B1 sky130_fd_sc_hd__buf_6
XFILLER_165_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_65_3 dadda_fa_3_65_3/A dadda_fa_3_65_3/B dadda_fa_3_65_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_66_1/B dadda_fa_4_65_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_58_2 dadda_fa_3_58_2/A dadda_fa_3_58_2/B dadda_fa_3_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_1/A dadda_fa_4_58_2/B sky130_fd_sc_hd__fa_1
XFILLER_120_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_28_0 dadda_fa_6_28_0/A dadda_fa_6_28_0/B dadda_fa_6_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_29_0/B dadda_fa_7_28_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_62_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2203 U$$2203/A U$$2253/B VGND VGND VPWR VPWR U$$2203/X sky130_fd_sc_hd__xor2_1
XU$$2214 U$$2625/A1 U$$2272/A2 U$$2625/B1 U$$2272/B2 VGND VGND VPWR VPWR U$$2215/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2225 U$$2225/A U$$2273/B VGND VGND VPWR VPWR U$$2225/X sky130_fd_sc_hd__xor2_1
XU$$2236 U$$44/A1 U$$2284/A2 U$$44/B1 U$$2284/B2 VGND VGND VPWR VPWR U$$2237/A sky130_fd_sc_hd__a22o_1
XU$$2247 U$$2247/A U$$2285/B VGND VGND VPWR VPWR U$$2247/X sky130_fd_sc_hd__xor2_1
XU$$1502 U$$2324/A1 U$$1502/A2 U$$1504/A1 U$$1502/B2 VGND VGND VPWR VPWR U$$1503/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2258 U$$888/A1 U$$2308/A2 U$$890/A1 U$$2308/B2 VGND VGND VPWR VPWR U$$2259/A sky130_fd_sc_hd__a22o_1
XU$$1513 U$$1513/A1 U$$1575/A2 U$$1515/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1514/A
+ sky130_fd_sc_hd__a22o_1
XU$$2269 U$$2269/A U$$2309/B VGND VGND VPWR VPWR U$$2269/X sky130_fd_sc_hd__xor2_1
XU$$1524 U$$1524/A U$$1558/B VGND VGND VPWR VPWR U$$1524/X sky130_fd_sc_hd__xor2_1
XFILLER_90_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1535 U$$987/A1 U$$1575/A2 U$$987/B1 U$$1575/B2 VGND VGND VPWR VPWR U$$1536/A sky130_fd_sc_hd__a22o_1
XFILLER_31_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1546 U$$1546/A U$$1546/B VGND VGND VPWR VPWR U$$1546/X sky130_fd_sc_hd__xor2_1
XFILLER_203_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1557 U$$461/A1 U$$1557/A2 U$$461/B1 U$$1557/B2 VGND VGND VPWR VPWR U$$1558/A sky130_fd_sc_hd__a22o_1
XFILLER_76_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1568 U$$1568/A U$$1592/B VGND VGND VPWR VPWR U$$1568/X sky130_fd_sc_hd__xor2_1
XU$$1579 U$$2949/A1 U$$1621/A2 U$$2951/A1 U$$1621/B2 VGND VGND VPWR VPWR U$$1580/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_229_ _358_/CLK _229_/D VGND VGND VPWR VPWR _229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_2 dadda_fa_2_60_2/A dadda_fa_2_60_2/B dadda_fa_2_60_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/A dadda_fa_3_60_3/A sky130_fd_sc_hd__fa_1
XFILLER_100_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater402 U$$689/X VGND VGND VPWR VPWR U$$793/A2 sky130_fd_sc_hd__buf_12
XFILLER_57_308 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$209 final_adder.U$$208/B final_adder.U$$979/B1 final_adder.U$$209/B1
+ VGND VGND VPWR VPWR final_adder.U$$209/X sky130_fd_sc_hd__a21o_1
Xrepeater413 U$$672/A2 VGND VGND VPWR VPWR U$$678/A2 sky130_fd_sc_hd__buf_12
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater424 U$$515/A2 VGND VGND VPWR VPWR U$$437/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_53_1 dadda_fa_2_53_1/A dadda_fa_2_53_1/B dadda_fa_2_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_0/CIN dadda_fa_3_53_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater435 U$$4238/A2 VGND VGND VPWR VPWR U$$4226/A2 sky130_fd_sc_hd__clkbuf_4
Xrepeater446 U$$4/X VGND VGND VPWR VPWR U$$94/A2 sky130_fd_sc_hd__buf_6
XFILLER_38_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater457 U$$3970/A2 VGND VGND VPWR VPWR U$$3874/A2 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_5_30_0 dadda_fa_5_30_0/A dadda_fa_5_30_0/B dadda_fa_5_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_31_0/A dadda_fa_6_30_0/CIN sky130_fd_sc_hd__fa_2
Xrepeater468 U$$3773/A2 VGND VGND VPWR VPWR U$$3739/A2 sky130_fd_sc_hd__buf_4
XU$$4150 input72/X U$$4188/A2 input73/X U$$4188/B2 VGND VGND VPWR VPWR U$$4151/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_46_0 U$$2759/X U$$2892/X U$$3025/X VGND VGND VPWR VPWR dadda_fa_3_47_0/B
+ dadda_fa_3_46_2/B sky130_fd_sc_hd__fa_1
Xrepeater479 U$$3429/X VGND VGND VPWR VPWR U$$3503/A2 sky130_fd_sc_hd__buf_4
XU$$4161 U$$4161/A U$$4243/B VGND VGND VPWR VPWR U$$4161/X sky130_fd_sc_hd__xor2_1
XFILLER_81_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4172 U$$4309/A1 U$$4176/A2 U$$4309/B1 U$$4176/B2 VGND VGND VPWR VPWR U$$4173/A
+ sky130_fd_sc_hd__a22o_1
XU$$4183 U$$4183/A U$$4227/B VGND VGND VPWR VPWR U$$4183/X sky130_fd_sc_hd__xor2_1
XFILLER_25_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4194 U$$4466/B1 U$$4210/A2 U$$4333/A1 U$$4210/B2 VGND VGND VPWR VPWR U$$4195/A
+ sky130_fd_sc_hd__a22o_1
XU$$3460 U$$3460/A U$$3480/B VGND VGND VPWR VPWR U$$3460/X sky130_fd_sc_hd__xor2_1
XU$$3471 U$$4430/A1 U$$3503/A2 U$$4432/A1 U$$3503/B2 VGND VGND VPWR VPWR U$$3472/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3482 U$$3482/A U$$3490/B VGND VGND VPWR VPWR U$$3482/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3493 U$$4176/B1 U$$3429/X U$$4178/B1 U$$3430/X VGND VGND VPWR VPWR U$$3494/A sky130_fd_sc_hd__a22o_1
XFILLER_34_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2770 U$$30/A1 U$$2782/A2 U$$32/A1 U$$2782/B2 VGND VGND VPWR VPWR U$$2771/A sky130_fd_sc_hd__a22o_1
XFILLER_22_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2781 U$$2781/A U$$2869/B VGND VGND VPWR VPWR U$$2781/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2792 U$$4297/B1 U$$2796/A2 U$$328/A1 U$$2796/B2 VGND VGND VPWR VPWR U$$2793/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_75_2 dadda_fa_4_75_2/A dadda_fa_4_75_2/B dadda_fa_4_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_76_0/CIN dadda_fa_5_75_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_68_1 dadda_fa_4_68_1/A dadda_fa_4_68_1/B dadda_fa_4_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/B dadda_fa_5_68_1/B sky130_fd_sc_hd__fa_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput205 c[53] VGND VGND VPWR VPWR input205/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_7_45_0 dadda_fa_7_45_0/A dadda_fa_7_45_0/B dadda_fa_7_45_0/CIN VGND VGND
+ VPWR VPWR _342_/D _213_/D sky130_fd_sc_hd__fa_2
Xinput216 c[63] VGND VGND VPWR VPWR input216/X sky130_fd_sc_hd__clkbuf_1
Xinput227 c[73] VGND VGND VPWR VPWR input227/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput238 c[83] VGND VGND VPWR VPWR input238/X sky130_fd_sc_hd__buf_2
XFILLER_76_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_1_35_0 U$$77/X U$$210/X VGND VGND VPWR VPWR dadda_fa_2_36_5/B dadda_fa_3_35_0/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$710 final_adder.U$$710/A final_adder.U$$710/B VGND VGND VPWR VPWR
+ final_adder.U$$790/A sky130_fd_sc_hd__and2_1
Xinput249 c[93] VGND VGND VPWR VPWR input249/X sky130_fd_sc_hd__clkbuf_4
XTAP_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$721 final_adder.U$$720/B final_adder.U$$617/X final_adder.U$$601/X
+ VGND VGND VPWR VPWR final_adder.U$$721/X sky130_fd_sc_hd__a21o_1
XTAP_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$743 final_adder.U$$742/B final_adder.U$$663/X final_adder.U$$631/X
+ VGND VGND VPWR VPWR final_adder.U$$743/X sky130_fd_sc_hd__a21o_1
XTAP_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$754 final_adder.U$$786/B final_adder.U$$754/B VGND VGND VPWR VPWR
+ final_adder.U$$754/X sky130_fd_sc_hd__and2_1
XFILLER_29_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$765 final_adder.U$$764/B final_adder.U$$685/X final_adder.U$$653/X
+ VGND VGND VPWR VPWR final_adder.U$$765/X sky130_fd_sc_hd__a21o_1
XFILLER_186_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$604 U$$56/A1 U$$636/A2 U$$878/B1 U$$636/B2 VGND VGND VPWR VPWR U$$605/A sky130_fd_sc_hd__a22o_1
XFILLER_90_108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$776 final_adder.U$$776/A final_adder.U$$776/B VGND VGND VPWR VPWR
+ final_adder.U$$776/X sky130_fd_sc_hd__and2_1
XU$$615 U$$615/A U$$617/B VGND VGND VPWR VPWR U$$615/X sky130_fd_sc_hd__xor2_1
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater980 U$$4045/A1 VGND VGND VPWR VPWR U$$4043/B1 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$787 final_adder.U$$786/B final_adder.U$$707/X final_adder.U$$675/X
+ VGND VGND VPWR VPWR final_adder.U$$787/X sky130_fd_sc_hd__a21o_1
Xrepeater991 input9/X VGND VGND VPWR VPWR U$$1209/B sky130_fd_sc_hd__buf_8
XU$$626 U$$763/A1 U$$672/A2 U$$763/B1 U$$668/B2 VGND VGND VPWR VPWR U$$627/A sky130_fd_sc_hd__a22o_1
XFILLER_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$798 final_adder.U$$798/A final_adder.U$$798/B VGND VGND VPWR VPWR
+ final_adder.U$$798/X sky130_fd_sc_hd__and2_1
XFILLER_71_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$637 U$$637/A U$$637/B VGND VGND VPWR VPWR U$$637/X sky130_fd_sc_hd__xor2_1
XU$$648 U$$783/B1 U$$652/A2 U$$650/A1 U$$652/B2 VGND VGND VPWR VPWR U$$649/A sky130_fd_sc_hd__a22o_1
XFILLER_72_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$659 U$$659/A U$$684/A VGND VGND VPWR VPWR U$$659/X sky130_fd_sc_hd__xor2_1
XFILLER_71_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_1188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1504 input123/X VGND VGND VPWR VPWR U$$3555/B1 sky130_fd_sc_hd__buf_4
XFILLER_158_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1515 U$$2318/B1 VGND VGND VPWR VPWR U$$950/A1 sky130_fd_sc_hd__buf_6
Xrepeater1526 U$$3852/B1 VGND VGND VPWR VPWR U$$4402/A1 sky130_fd_sc_hd__buf_6
Xrepeater1537 U$$136/A VGND VGND VPWR VPWR U$$3/A sky130_fd_sc_hd__buf_4
XFILLER_126_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1548 U$$2316/A1 VGND VGND VPWR VPWR U$$946/A1 sky130_fd_sc_hd__buf_6
Xrepeater1559 U$$1764/B1 VGND VGND VPWR VPWR U$$2312/B1 sky130_fd_sc_hd__buf_6
XFILLER_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_70_1 dadda_fa_3_70_1/A dadda_fa_3_70_1/B dadda_fa_3_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_0/CIN dadda_fa_4_70_2/A sky130_fd_sc_hd__fa_1
XFILLER_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_63_0 dadda_fa_3_63_0/A dadda_fa_3_63_0/B dadda_fa_3_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_0/B dadda_fa_4_63_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2000 U$$2409/B1 U$$2040/A2 U$$3235/A1 U$$2040/B2 VGND VGND VPWR VPWR U$$2001/A
+ sky130_fd_sc_hd__a22o_1
XU$$2011 U$$2011/A U$$2037/B VGND VGND VPWR VPWR U$$2011/X sky130_fd_sc_hd__xor2_1
XFILLER_165_1206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2022 U$$789/A1 U$$2022/A2 U$$928/A1 U$$2022/B2 VGND VGND VPWR VPWR U$$2023/A sky130_fd_sc_hd__a22o_1
XFILLER_62_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2033 U$$2033/A U$$2047/B VGND VGND VPWR VPWR U$$2033/X sky130_fd_sc_hd__xor2_1
XFILLER_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2044 U$$948/A1 U$$1922/X U$$2044/B1 U$$1923/X VGND VGND VPWR VPWR U$$2045/A sky130_fd_sc_hd__a22o_1
XU$$1310 U$$1310/A U$$1316/B VGND VGND VPWR VPWR U$$1310/X sky130_fd_sc_hd__xor2_1
XU$$2055 input22/X VGND VGND VPWR VPWR U$$2055/Y sky130_fd_sc_hd__inv_1
XFILLER_74_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1321 U$$2415/B1 U$$1353/A2 U$$2282/A1 U$$1349/B2 VGND VGND VPWR VPWR U$$1322/A
+ sky130_fd_sc_hd__a22o_1
XU$$2066 U$$2066/A U$$2094/B VGND VGND VPWR VPWR U$$2066/X sky130_fd_sc_hd__xor2_1
XU$$1332 U$$1332/A U$$1338/B VGND VGND VPWR VPWR U$$1332/X sky130_fd_sc_hd__xor2_1
XU$$2077 U$$2625/A1 U$$2093/A2 U$$2625/B1 U$$2093/B2 VGND VGND VPWR VPWR U$$2078/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2088 U$$2088/A U$$2092/B VGND VGND VPWR VPWR U$$2088/X sky130_fd_sc_hd__xor2_1
XFILLER_50_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1343 U$$932/A1 U$$1353/A2 U$$932/B1 U$$1238/X VGND VGND VPWR VPWR U$$1344/A sky130_fd_sc_hd__a22o_1
XFILLER_200_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1354 U$$1354/A U$$1354/B VGND VGND VPWR VPWR U$$1354/X sky130_fd_sc_hd__xor2_1
XFILLER_210_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2099 U$$3878/B1 U$$2099/A2 U$$44/B1 U$$2099/B2 VGND VGND VPWR VPWR U$$2100/A sky130_fd_sc_hd__a22o_1
XFILLER_128_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1365 U$$2324/A1 U$$1367/A2 U$$1504/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1366/A
+ sky130_fd_sc_hd__a22o_1
XU$$1376 U$$1376/A1 U$$1404/A2 U$$1515/A1 U$$1404/B2 VGND VGND VPWR VPWR U$$1377/A
+ sky130_fd_sc_hd__a22o_1
XU$$1387 U$$1387/A U$$1399/B VGND VGND VPWR VPWR U$$1387/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_120_0 dadda_fa_7_120_0/A dadda_fa_7_120_0/B dadda_fa_7_120_0/CIN VGND
+ VGND VPWR VPWR _417_/D _288_/D sky130_fd_sc_hd__fa_1
XU$$1398 U$$987/A1 U$$1404/A2 U$$987/B1 U$$1404/B2 VGND VGND VPWR VPWR U$$1399/A sky130_fd_sc_hd__a22o_1
XFILLER_88_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_85_1 dadda_fa_5_85_1/A dadda_fa_5_85_1/B dadda_fa_5_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_86_0/B dadda_fa_7_85_0/A sky130_fd_sc_hd__fa_1
XFILLER_102_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_78_0 dadda_fa_5_78_0/A dadda_fa_5_78_0/B dadda_fa_5_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_79_0/A dadda_fa_6_78_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_144_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_77_8 input231/X dadda_fa_1_77_8/B dadda_fa_1_77_8/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_78_3/A dadda_fa_3_77_0/A sky130_fd_sc_hd__fa_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$50 _346_/Q _218_/Q VGND VGND VPWR VPWR final_adder.U$$975/B1 final_adder.U$$204/A
+ sky130_fd_sc_hd__ha_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$61 _357_/Q _229_/Q VGND VGND VPWR VPWR final_adder.U$$195/B1 final_adder.U$$194/B
+ sky130_fd_sc_hd__ha_1
XFILLER_80_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3290 input44/X VGND VGND VPWR VPWR U$$3290/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$72 _368_/Q _240_/Q VGND VGND VPWR VPWR final_adder.U$$953/B1 final_adder.U$$182/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$83 _379_/Q _251_/Q VGND VGND VPWR VPWR final_adder.U$$173/B1 final_adder.U$$172/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$94 _390_/Q _262_/Q VGND VGND VPWR VPWR final_adder.U$$931/B1 final_adder.U$$160/A
+ sky130_fd_sc_hd__ha_1
XFILLER_80_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1650_1721 VGND VGND VPWR VPWR U$$1650_1721/HI U$$1650/A1 sky130_fd_sc_hd__conb_1
XFILLER_108_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_80_0 dadda_fa_4_80_0/A dadda_fa_4_80_0/B dadda_fa_4_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/A dadda_fa_5_80_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_101_3 dadda_fa_3_101_3/A dadda_fa_3_101_3/B dadda_fa_3_101_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_102_1/B dadda_fa_4_101_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_87 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_20 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$540 final_adder.U$$548/B final_adder.U$$540/B VGND VGND VPWR VPWR
+ final_adder.U$$660/B sky130_fd_sc_hd__and2_1
XTAP_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$551 final_adder.U$$550/B final_adder.U$$435/X final_adder.U$$427/X
+ VGND VGND VPWR VPWR final_adder.U$$551/X sky130_fd_sc_hd__a21o_1
XTAP_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$562 final_adder.U$$570/B final_adder.U$$562/B VGND VGND VPWR VPWR
+ final_adder.U$$682/B sky130_fd_sc_hd__and2_1
Xdadda_fa_6_108_0 dadda_fa_6_108_0/A dadda_fa_6_108_0/B dadda_fa_6_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_109_0/B dadda_fa_7_108_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$401 U$$401/A U$$411/A VGND VGND VPWR VPWR U$$401/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$573 final_adder.U$$572/B final_adder.U$$457/X final_adder.U$$449/X
+ VGND VGND VPWR VPWR final_adder.U$$573/X sky130_fd_sc_hd__a21o_1
XTAP_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$412 U$$412/A VGND VGND VPWR VPWR U$$414/B sky130_fd_sc_hd__inv_1
XFILLER_45_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$584 final_adder.U$$592/B final_adder.U$$584/B VGND VGND VPWR VPWR
+ final_adder.U$$704/B sky130_fd_sc_hd__and2_1
XU$$423 U$$969/B1 U$$437/A2 U$$836/A1 U$$437/B2 VGND VGND VPWR VPWR U$$424/A sky130_fd_sc_hd__a22o_1
XTAP_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$595 final_adder.U$$594/B final_adder.U$$479/X final_adder.U$$471/X
+ VGND VGND VPWR VPWR final_adder.U$$595/X sky130_fd_sc_hd__a21o_1
XU$$434 U$$434/A U$$436/B VGND VGND VPWR VPWR U$$434/X sky130_fd_sc_hd__xor2_1
XTAP_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$445 U$$34/A1 U$$515/A2 U$$36/A1 U$$515/B2 VGND VGND VPWR VPWR U$$446/A sky130_fd_sc_hd__a22o_1
XTAP_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$456 U$$456/A U$$492/B VGND VGND VPWR VPWR U$$456/X sky130_fd_sc_hd__xor2_1
XFILLER_205_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_28_3 dadda_fa_3_28_3/A dadda_fa_3_28_3/B dadda_fa_3_28_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_29_1/B dadda_fa_4_28_2/CIN sky130_fd_sc_hd__fa_1
XU$$467 U$$56/A1 U$$483/A2 U$$878/B1 U$$483/B2 VGND VGND VPWR VPWR U$$468/A sky130_fd_sc_hd__a22o_1
XFILLER_71_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$478 U$$478/A U$$504/B VGND VGND VPWR VPWR U$$478/X sky130_fd_sc_hd__xor2_1
XU$$489 U$$763/A1 U$$491/A2 U$$763/B1 U$$491/B2 VGND VGND VPWR VPWR U$$490/A sky130_fd_sc_hd__a22o_1
XFILLER_185_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_371 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_95_0 dadda_fa_6_95_0/A dadda_fa_6_95_0/B dadda_fa_6_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_96_0/B dadda_fa_7_95_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_139_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_994 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1301 U$$3510/B VGND VGND VPWR VPWR U$$3518/B sky130_fd_sc_hd__buf_12
XFILLER_201_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1312 U$$3228/B VGND VGND VPWR VPWR U$$3188/B sky130_fd_sc_hd__buf_6
XFILLER_201_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1323 U$$3109/B VGND VGND VPWR VPWR U$$3077/B sky130_fd_sc_hd__buf_12
Xrepeater1334 U$$2978/B VGND VGND VPWR VPWR U$$2968/B sky130_fd_sc_hd__buf_12
XFILLER_158_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1345 U$$2876/A VGND VGND VPWR VPWR U$$2859/B sky130_fd_sc_hd__buf_6
XFILLER_10_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1356 U$$272/B VGND VGND VPWR VPWR U$$264/B sky130_fd_sc_hd__buf_8
XFILLER_113_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1367 U$$2602/A VGND VGND VPWR VPWR U$$2601/B sky130_fd_sc_hd__buf_8
XFILLER_119_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1378 U$$821/A VGND VGND VPWR VPWR U$$794/B sky130_fd_sc_hd__buf_12
XFILLER_125_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1389 U$$2465/A VGND VGND VPWR VPWR U$$2380/B sky130_fd_sc_hd__buf_8
XFILLER_107_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_30_3 U$$1264/X U$$1397/X U$$1530/X VGND VGND VPWR VPWR dadda_fa_3_31_2/A
+ dadda_fa_3_30_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_165_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$990 U$$990/A U$$994/B VGND VGND VPWR VPWR U$$990/X sky130_fd_sc_hd__xor2_1
XFILLER_211_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1140 U$$44/A1 U$$1174/A2 U$$46/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1141/A sky130_fd_sc_hd__a22o_1
XFILLER_211_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1151 U$$1151/A U$$1195/B VGND VGND VPWR VPWR U$$1151/X sky130_fd_sc_hd__xor2_1
XFILLER_50_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1162 U$$888/A1 U$$1162/A2 U$$890/A1 U$$1162/B2 VGND VGND VPWR VPWR U$$1163/A sky130_fd_sc_hd__a22o_1
XU$$1173 U$$1173/A U$$1175/B VGND VGND VPWR VPWR U$$1173/X sky130_fd_sc_hd__xor2_1
XFILLER_149_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1184 U$$3922/B1 U$$1222/A2 U$$3787/B1 U$$1222/B2 VGND VGND VPWR VPWR U$$1185/A
+ sky130_fd_sc_hd__a22o_1
XU$$1195 U$$1195/A U$$1195/B VGND VGND VPWR VPWR U$$1195/X sky130_fd_sc_hd__xor2_1
XFILLER_31_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_82_6 U$$3629/X U$$3762/X U$$3895/X VGND VGND VPWR VPWR dadda_fa_2_83_3/B
+ dadda_fa_2_82_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_75_5 U$$3615/X U$$3748/X U$$3881/X VGND VGND VPWR VPWR dadda_fa_2_76_2/A
+ dadda_fa_2_75_5/A sky130_fd_sc_hd__fa_1
XFILLER_86_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_723 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_4 U$$4133/X U$$4266/X U$$4399/X VGND VGND VPWR VPWR dadda_fa_2_69_1/CIN
+ dadda_fa_2_68_4/CIN sky130_fd_sc_hd__fa_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_38_2 dadda_fa_4_38_2/A dadda_fa_4_38_2/B dadda_fa_4_38_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_39_0/CIN dadda_fa_5_38_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 _384_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _366_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_1103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_923 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_476 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_3 U$$1330/X U$$1463/X U$$1596/X VGND VGND VPWR VPWR dadda_fa_1_64_6/B
+ dadda_fa_1_63_8/B sky130_fd_sc_hd__fa_1
XTAP_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_40_2 dadda_fa_3_40_2/A dadda_fa_3_40_2/B dadda_fa_3_40_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_1/A dadda_fa_4_40_2/B sky130_fd_sc_hd__fa_1
XTAP_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$370 final_adder.U$$372/B final_adder.U$$370/B VGND VGND VPWR VPWR
+ final_adder.U$$496/B sky130_fd_sc_hd__and2_1
XTAP_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$381 final_adder.U$$378/A final_adder.U$$255/X final_adder.U$$253/X
+ VGND VGND VPWR VPWR final_adder.U$$381/X sky130_fd_sc_hd__a21o_2
XTAP_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$220 U$$220/A U$$264/B VGND VGND VPWR VPWR U$$220/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_33_1 dadda_fa_3_33_1/A dadda_fa_3_33_1/B dadda_fa_3_33_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_0/CIN dadda_fa_4_33_2/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$392 final_adder.U$$396/B final_adder.U$$392/B VGND VGND VPWR VPWR
+ final_adder.U$$516/B sky130_fd_sc_hd__and2_1
XTAP_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$231 U$$94/A1 U$$263/A2 U$$96/A1 U$$231/B2 VGND VGND VPWR VPWR U$$232/A sky130_fd_sc_hd__a22o_1
XFILLER_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$242 U$$242/A U$$244/B VGND VGND VPWR VPWR U$$242/X sky130_fd_sc_hd__xor2_1
XFILLER_45_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_10_0 dadda_fa_6_10_0/A dadda_fa_6_10_0/B dadda_fa_6_10_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_11_0/B dadda_fa_7_10_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$253 U$$388/B1 U$$257/A2 U$$392/A1 U$$257/B2 VGND VGND VPWR VPWR U$$254/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_26_0 U$$1123/X U$$1256/X U$$1389/X VGND VGND VPWR VPWR dadda_fa_4_27_0/B
+ dadda_fa_4_26_1/CIN sky130_fd_sc_hd__fa_1
XTAP_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$264 U$$264/A U$$264/B VGND VGND VPWR VPWR U$$264/X sky130_fd_sc_hd__xor2_1
XFILLER_75_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$275 U$$275/A VGND VGND VPWR VPWR U$$277/B sky130_fd_sc_hd__inv_1
XFILLER_72_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$286 U$$12/A1 U$$316/A2 U$$14/A1 U$$316/B2 VGND VGND VPWR VPWR U$$287/A sky130_fd_sc_hd__a22o_1
XFILLER_44_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$297 U$$297/A U$$379/B VGND VGND VPWR VPWR U$$297/X sky130_fd_sc_hd__xor2_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_583 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_931 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3 U$$3/A U$$3/B VGND VGND VPWR VPWR U$$3/X sky130_fd_sc_hd__and2_1
XFILLER_127_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput306 output306/A VGND VGND VPWR VPWR o[29] sky130_fd_sc_hd__buf_2
Xdadda_fa_2_92_5 dadda_fa_2_92_5/A dadda_fa_2_92_5/B dadda_fa_2_92_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_93_2/A dadda_fa_4_92_0/A sky130_fd_sc_hd__fa_1
Xrepeater1120 input74/X VGND VGND VPWR VPWR U$$4015/B1 sky130_fd_sc_hd__buf_6
Xoutput317 output317/A VGND VGND VPWR VPWR o[39] sky130_fd_sc_hd__buf_2
Xrepeater1131 U$$38/B1 VGND VGND VPWR VPWR U$$40/A1 sky130_fd_sc_hd__buf_4
Xoutput328 output328/A VGND VGND VPWR VPWR o[49] sky130_fd_sc_hd__buf_2
XU$$4471_1812 VGND VGND VPWR VPWR U$$4471_1812/HI U$$4471/B sky130_fd_sc_hd__conb_1
Xrepeater1142 U$$4422/A1 VGND VGND VPWR VPWR U$$4011/A1 sky130_fd_sc_hd__buf_6
XFILLER_114_614 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1153 input70/X VGND VGND VPWR VPWR U$$4146/A1 sky130_fd_sc_hd__clkbuf_8
Xoutput339 output339/A VGND VGND VPWR VPWR o[59] sky130_fd_sc_hd__buf_2
XFILLER_141_411 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_85_4 dadda_fa_2_85_4/A dadda_fa_2_85_4/B dadda_fa_2_85_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_1/CIN dadda_fa_3_85_3/CIN sky130_fd_sc_hd__fa_1
Xrepeater1164 U$$3183/B1 VGND VGND VPWR VPWR U$$854/B1 sky130_fd_sc_hd__buf_4
XFILLER_153_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1175 U$$4005/A1 VGND VGND VPWR VPWR U$$3183/A1 sky130_fd_sc_hd__buf_6
XFILLER_113_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1186 U$$4275/B1 VGND VGND VPWR VPWR U$$3727/B1 sky130_fd_sc_hd__buf_8
Xrepeater1197 U$$967/A1 VGND VGND VPWR VPWR U$$8/A1 sky130_fd_sc_hd__buf_2
XFILLER_4_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_78_3 dadda_fa_2_78_3/A dadda_fa_2_78_3/B dadda_fa_2_78_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/B dadda_fa_3_78_3/B sky130_fd_sc_hd__fa_1
XFILLER_45_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_48_1 dadda_fa_5_48_1/A dadda_fa_5_48_1/B dadda_fa_5_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_49_0/B dadda_fa_7_48_0/A sky130_fd_sc_hd__fa_1
XFILLER_83_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_992 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3970_1756 VGND VGND VPWR VPWR U$$3970_1756/HI U$$3970/B1 sky130_fd_sc_hd__conb_1
XFILLER_36_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_101_2 U$$3401/X U$$3534/X U$$3667/X VGND VGND VPWR VPWR dadda_fa_3_102_2/B
+ dadda_fa_3_101_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_1041 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_122_1 input154/X dadda_fa_5_122_1/B dadda_ha_4_122_0/SUM VGND VGND VPWR
+ VPWR dadda_fa_6_123_0/B dadda_fa_7_122_0/A sky130_fd_sc_hd__fa_1
XFILLER_177_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_115_0 dadda_fa_5_115_0/A dadda_fa_5_115_0/B dadda_fa_5_115_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_116_0/A dadda_fa_6_115_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_80_3 U$$2295/X U$$2428/X U$$2561/X VGND VGND VPWR VPWR dadda_fa_2_81_1/CIN
+ dadda_fa_2_80_4/B sky130_fd_sc_hd__fa_1
XFILLER_160_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_73_2 U$$2680/X U$$2813/X U$$2946/X VGND VGND VPWR VPWR dadda_fa_2_74_1/A
+ dadda_fa_2_73_4/A sky130_fd_sc_hd__fa_1
XFILLER_58_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_50_1 dadda_fa_4_50_1/A dadda_fa_4_50_1/B dadda_fa_4_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/B dadda_fa_5_50_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_66_1 U$$2932/X U$$3065/X U$$3198/X VGND VGND VPWR VPWR dadda_fa_2_67_0/CIN
+ dadda_fa_2_66_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_ha_2_100_4 U$$4064/X U$$4197/X VGND VGND VPWR VPWR dadda_fa_3_101_2/CIN dadda_fa_4_100_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_24_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_43_0 dadda_fa_4_43_0/A dadda_fa_4_43_0/B dadda_fa_4_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/A dadda_fa_5_43_1/A sky130_fd_sc_hd__fa_1
XFILLER_101_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_59_0 U$$1588/X U$$1721/X U$$1854/X VGND VGND VPWR VPWR dadda_fa_2_60_0/B
+ dadda_fa_2_59_3/B sky130_fd_sc_hd__fa_1
XFILLER_101_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_400_ _401_/CLK _400_/D VGND VGND VPWR VPWR _400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1909 U$$2044/B1 U$$1785/X U$$4514/A1 U$$1786/X VGND VGND VPWR VPWR U$$1910/A sky130_fd_sc_hd__a22o_1
XFILLER_42_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_859 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_331_ _337_/CLK _331_/D VGND VGND VPWR VPWR _331_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1048 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_262_ _407_/CLK _262_/D VGND VGND VPWR VPWR _262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_391 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_193_ _323_/CLK _193_/D VGND VGND VPWR VPWR _193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_95_3 dadda_fa_3_95_3/A dadda_fa_3_95_3/B dadda_fa_3_95_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_96_1/B dadda_fa_4_95_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_88_2 dadda_fa_3_88_2/A dadda_fa_3_88_2/B dadda_fa_3_88_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_1/A dadda_fa_4_88_2/B sky130_fd_sc_hd__fa_1
XFILLER_124_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_0_55_1 U$$516/X U$$649/X VGND VGND VPWR VPWR dadda_fa_1_56_8/A dadda_fa_2_55_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_58_0 dadda_fa_6_58_0/A dadda_fa_6_58_0/B dadda_fa_6_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_59_0/B dadda_fa_7_58_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater809 U$$2302/B2 VGND VGND VPWR VPWR U$$2272/B2 sky130_fd_sc_hd__buf_6
XU$$4502 U$$4502/A1 U$$4388/X U$$4504/A1 U$$4512/B2 VGND VGND VPWR VPWR U$$4503/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4513 U$$4513/A U$$4513/B VGND VGND VPWR VPWR U$$4513/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_61_0 U$$129/X U$$262/X U$$395/X VGND VGND VPWR VPWR dadda_fa_1_62_5/CIN
+ dadda_fa_1_61_7/CIN sky130_fd_sc_hd__fa_1
XU$$3801 U$$4210/B1 U$$3813/A2 U$$3801/B1 U$$3813/B2 VGND VGND VPWR VPWR U$$3802/A
+ sky130_fd_sc_hd__a22o_1
XU$$16 U$$16/A1 U$$8/A2 U$$18/A1 U$$8/B2 VGND VGND VPWR VPWR U$$17/A sky130_fd_sc_hd__a22o_1
XFILLER_65_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3812 U$$3812/A U$$3814/B VGND VGND VPWR VPWR U$$3812/X sky130_fd_sc_hd__xor2_1
XTAP_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$27 U$$27/A U$$43/B VGND VGND VPWR VPWR U$$27/X sky130_fd_sc_hd__xor2_1
XTAP_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3823 U$$3960/A1 U$$3833/A2 U$$3960/B1 U$$3833/B2 VGND VGND VPWR VPWR U$$3824/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_117_2 U$$4497/X input148/X dadda_fa_4_117_2/CIN VGND VGND VPWR VPWR dadda_fa_5_118_0/CIN
+ dadda_fa_5_117_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$38 U$$38/A1 U$$42/A2 U$$38/B1 U$$42/B2 VGND VGND VPWR VPWR U$$39/A sky130_fd_sc_hd__a22o_1
XFILLER_65_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3834 U$$3834/A U$$3834/B VGND VGND VPWR VPWR U$$3834/X sky130_fd_sc_hd__xor2_1
XU$$49 U$$49/A U$$51/B VGND VGND VPWR VPWR U$$49/X sky130_fd_sc_hd__xor2_1
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3845 U$$3845/A U$$3879/B VGND VGND VPWR VPWR U$$3845/X sky130_fd_sc_hd__xor2_1
XTAP_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3856 U$$4402/B1 U$$3874/A2 U$$4269/A1 U$$3874/B2 VGND VGND VPWR VPWR U$$3857/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3867 U$$3867/A U$$3903/B VGND VGND VPWR VPWR U$$3867/X sky130_fd_sc_hd__xor2_1
XTAP_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3878 U$$4289/A1 U$$3878/A2 U$$3878/B1 U$$3878/B2 VGND VGND VPWR VPWR U$$3879/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3889 U$$3889/A U$$3971/B VGND VGND VPWR VPWR U$$3889/X sky130_fd_sc_hd__xor2_1
XFILLER_127_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4429_1791 VGND VGND VPWR VPWR U$$4429_1791/HI U$$4429/B sky130_fd_sc_hd__conb_1
XFILLER_127_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_18 _332_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _338_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_203_1025 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_90_2 U$$4044/X U$$4177/X U$$4310/X VGND VGND VPWR VPWR dadda_fa_3_91_1/A
+ dadda_fa_3_90_3/A sky130_fd_sc_hd__fa_1
XFILLER_177_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_83_1 input238/X dadda_fa_2_83_1/B dadda_fa_2_83_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_84_0/CIN dadda_fa_3_83_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_142_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_60_0 dadda_fa_5_60_0/A dadda_fa_5_60_0/B dadda_fa_5_60_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_61_0/A dadda_fa_6_60_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_76_0 dadda_fa_2_76_0/A dadda_fa_2_76_0/B dadda_fa_2_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_0/B dadda_fa_3_76_2/B sky130_fd_sc_hd__fa_1
XFILLER_102_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_52_7 U$$3170/X U$$3303/X U$$3436/X VGND VGND VPWR VPWR dadda_fa_2_53_2/CIN
+ dadda_fa_2_52_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2883_1741 VGND VGND VPWR VPWR U$$2883_1741/HI U$$2883/A1 sky130_fd_sc_hd__conb_1
XFILLER_55_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_1231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_98_1 dadda_fa_4_98_1/A dadda_fa_4_98_1/B dadda_fa_4_98_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/B dadda_fa_5_98_1/B sky130_fd_sc_hd__fa_1
XFILLER_192_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_75_0 dadda_fa_7_75_0/A dadda_fa_7_75_0/B dadda_fa_7_75_0/CIN VGND VGND
+ VPWR VPWR _372_/D _243_/D sky130_fd_sc_hd__fa_1
XFILLER_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3108 U$$3108/A1 U$$3108/A2 U$$3108/B1 U$$3108/B2 VGND VGND VPWR VPWR U$$3109/A
+ sky130_fd_sc_hd__a22o_1
XU$$3119 U$$3119/A U$$3133/B VGND VGND VPWR VPWR U$$3119/X sky130_fd_sc_hd__xor2_1
XFILLER_207_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2407 U$$2955/A1 U$$2435/A2 U$$3366/B1 U$$2435/B2 VGND VGND VPWR VPWR U$$2408/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2418 U$$2418/A U$$2426/B VGND VGND VPWR VPWR U$$2418/X sky130_fd_sc_hd__xor2_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2429 U$$3114/A1 U$$2449/A2 U$$3116/A1 U$$2449/B2 VGND VGND VPWR VPWR U$$2430/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1706 U$$3348/B1 U$$1706/A2 U$$3215/A1 U$$1706/B2 VGND VGND VPWR VPWR U$$1707/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1717 U$$1717/A U$$1765/B VGND VGND VPWR VPWR U$$1717/X sky130_fd_sc_hd__xor2_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1728 U$$630/B1 U$$1736/A2 U$$86/A1 U$$1736/B2 VGND VGND VPWR VPWR U$$1729/A sky130_fd_sc_hd__a22o_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1739 U$$1739/A U$$1739/B VGND VGND VPWR VPWR U$$1739/X sky130_fd_sc_hd__xor2_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_314_ _314_/CLK _314_/D VGND VGND VPWR VPWR _314_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_245_ _376_/CLK _245_/D VGND VGND VPWR VPWR _245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput16 a[23] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput27 a[33] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__buf_6
XFILLER_195_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 a[43] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__buf_6
X_176_ _326_/CLK _176_/D VGND VGND VPWR VPWR _176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput49 a[53] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__buf_6
XFILLER_196_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_93_0 dadda_fa_3_93_0/A dadda_fa_3_93_0/B dadda_fa_3_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_0/B dadda_fa_4_93_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_202_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_786 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater606 U$$1511/X VGND VGND VPWR VPWR U$$1607/A2 sky130_fd_sc_hd__buf_6
XFILLER_96_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater617 U$$1504/A2 VGND VGND VPWR VPWR U$$1502/A2 sky130_fd_sc_hd__buf_6
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater628 U$$1337/A2 VGND VGND VPWR VPWR U$$1289/A2 sky130_fd_sc_hd__buf_4
XU$$4310 U$$4310/A U$$4310/B VGND VGND VPWR VPWR U$$4310/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_55_5 dadda_fa_2_55_5/A dadda_fa_2_55_5/B dadda_fa_2_55_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_56_2/A dadda_fa_4_55_0/A sky130_fd_sc_hd__fa_1
XU$$4321 U$$4458/A1 U$$4327/A2 U$$4460/A1 U$$4327/B2 VGND VGND VPWR VPWR U$$4322/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater639 U$$1100/X VGND VGND VPWR VPWR U$$1204/A2 sky130_fd_sc_hd__buf_8
XFILLER_120_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4332 U$$4332/A U$$4354/B VGND VGND VPWR VPWR U$$4332/X sky130_fd_sc_hd__xor2_1
XU$$4343 U$$4343/A1 U$$4349/A2 U$$4343/B1 U$$4349/B2 VGND VGND VPWR VPWR U$$4344/A
+ sky130_fd_sc_hd__a22o_1
XU$$4354 U$$4354/A U$$4354/B VGND VGND VPWR VPWR U$$4354/X sky130_fd_sc_hd__xor2_1
XU$$4365 U$$4502/A1 U$$4369/A2 U$$4365/B1 U$$4369/B2 VGND VGND VPWR VPWR U$$4366/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_48_4 dadda_fa_2_48_4/A dadda_fa_2_48_4/B dadda_fa_2_48_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_1/CIN dadda_fa_3_48_3/CIN sky130_fd_sc_hd__fa_1
XU$$3620 input82/X U$$3644/A2 input83/X U$$3644/B2 VGND VGND VPWR VPWR U$$3621/A sky130_fd_sc_hd__a22o_1
XU$$3631 U$$3631/A U$$3637/B VGND VGND VPWR VPWR U$$3631/X sky130_fd_sc_hd__xor2_1
XFILLER_77_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4376 U$$4376/A U$$4382/B VGND VGND VPWR VPWR U$$4376/X sky130_fd_sc_hd__xor2_1
XFILLER_92_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4387 U$$4387/A U$$4387/B VGND VGND VPWR VPWR U$$4387/X sky130_fd_sc_hd__and2_1
XU$$3642 U$$3642/A1 U$$3566/X U$$3644/A1 U$$3567/X VGND VGND VPWR VPWR U$$3643/A sky130_fd_sc_hd__a22o_1
XU$$3653 U$$3653/A U$$3683/B VGND VGND VPWR VPWR U$$3653/X sky130_fd_sc_hd__xor2_1
XU$$4398 U$$4398/A1 U$$4388/X U$$4400/A1 U$$4432/B2 VGND VGND VPWR VPWR U$$4399/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3664 U$$4210/B1 U$$3680/A2 U$$3801/B1 U$$3680/B2 VGND VGND VPWR VPWR U$$3665/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3675 U$$3675/A U$$3683/B VGND VGND VPWR VPWR U$$3675/X sky130_fd_sc_hd__xor2_1
XU$$2930 U$$2930/A U$$2968/B VGND VGND VPWR VPWR U$$2930/X sky130_fd_sc_hd__xor2_1
XFILLER_46_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3686 input118/X U$$3686/A2 input119/X U$$3686/B2 VGND VGND VPWR VPWR U$$3687/A
+ sky130_fd_sc_hd__a22o_1
XU$$2941 U$$3213/B1 U$$2949/A2 U$$4450/A1 U$$2949/B2 VGND VGND VPWR VPWR U$$2942/A
+ sky130_fd_sc_hd__a22o_1
XU$$3697 U$$3697/A U$$3697/B VGND VGND VPWR VPWR U$$3697/X sky130_fd_sc_hd__xor2_1
XU$$2952 U$$2952/A U$$2996/B VGND VGND VPWR VPWR U$$2952/X sky130_fd_sc_hd__xor2_1
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2963 U$$3511/A1 U$$2985/A2 U$$3648/B1 U$$2882/X VGND VGND VPWR VPWR U$$2964/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2974 U$$2974/A U$$2978/B VGND VGND VPWR VPWR U$$2974/X sky130_fd_sc_hd__xor2_1
XU$$2985 U$$517/B1 U$$2985/A2 U$$384/A1 U$$2985/B2 VGND VGND VPWR VPWR U$$2986/A sky130_fd_sc_hd__a22o_1
XU$$2996 U$$2996/A U$$2996/B VGND VGND VPWR VPWR U$$2996/X sky130_fd_sc_hd__xor2_1
XFILLER_166_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_915 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_1_44_5 U$$2090/X U$$2223/X VGND VGND VPWR VPWR dadda_fa_2_45_4/A dadda_fa_3_44_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_25_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$903 final_adder.U$$132/A final_adder.U$$841/X final_adder.U$$903/B1
+ VGND VGND VPWR VPWR final_adder.U$$903/X sky130_fd_sc_hd__a21o_1
XTAP_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$925 final_adder.U$$154/A final_adder.U$$863/X final_adder.U$$925/B1
+ VGND VGND VPWR VPWR final_adder.U$$925/X sky130_fd_sc_hd__a21o_1
XFILLER_68_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$947 final_adder.U$$176/A final_adder.U$$885/X final_adder.U$$947/B1
+ VGND VGND VPWR VPWR final_adder.U$$947/X sky130_fd_sc_hd__a21o_1
XFILLER_21_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_50_4 U$$1703/X U$$1836/X U$$1969/X VGND VGND VPWR VPWR dadda_fa_2_51_1/CIN
+ dadda_fa_2_50_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$808 U$$808/A U$$808/B VGND VGND VPWR VPWR U$$808/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$969 final_adder.U$$198/A final_adder.U$$811/X final_adder.U$$969/B1
+ VGND VGND VPWR VPWR final_adder.U$$969/X sky130_fd_sc_hd__a21o_1
XU$$819 U$$956/A1 U$$689/X U$$819/B1 U$$690/X VGND VGND VPWR VPWR U$$820/A sky130_fd_sc_hd__a22o_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_43_3 U$$1290/X U$$1423/X U$$1556/X VGND VGND VPWR VPWR dadda_fa_2_44_3/CIN
+ dadda_fa_2_43_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_20_2 dadda_fa_4_20_2/A dadda_fa_4_20_2/B dadda_ha_3_20_3/SUM VGND VGND
+ VPWR VPWR dadda_fa_5_21_0/CIN dadda_fa_5_20_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_189_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_13_1 U$$432/X U$$565/X U$$698/X VGND VGND VPWR VPWR dadda_fa_5_14_0/B
+ dadda_fa_5_13_1/B sky130_fd_sc_hd__fa_1
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_1023 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1708 input100/X VGND VGND VPWR VPWR U$$4335/B1 sky130_fd_sc_hd__buf_6
XFILLER_164_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1046 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_607 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_58_3 dadda_fa_3_58_3/A dadda_fa_3_58_3/B dadda_fa_3_58_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_59_1/B dadda_fa_4_58_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2204 U$$3300/A1 U$$2252/A2 U$$3300/B1 U$$2252/B2 VGND VGND VPWR VPWR U$$2205/A
+ sky130_fd_sc_hd__a22o_1
XU$$2215 U$$2215/A U$$2273/B VGND VGND VPWR VPWR U$$2215/X sky130_fd_sc_hd__xor2_1
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2226 U$$4144/A1 U$$2226/A2 U$$4144/B1 U$$2226/B2 VGND VGND VPWR VPWR U$$2227/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2237 U$$2237/A U$$2285/B VGND VGND VPWR VPWR U$$2237/X sky130_fd_sc_hd__xor2_1
XU$$1503 U$$1503/A U$$1507/A VGND VGND VPWR VPWR U$$1503/X sky130_fd_sc_hd__xor2_1
XU$$2248 input81/X U$$2284/A2 U$$3618/B1 U$$2284/B2 VGND VGND VPWR VPWR U$$2249/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2259 U$$2259/A U$$2309/B VGND VGND VPWR VPWR U$$2259/X sky130_fd_sc_hd__xor2_1
XFILLER_76_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1514 U$$1514/A U$$1574/B VGND VGND VPWR VPWR U$$1514/X sky130_fd_sc_hd__xor2_1
XU$$1525 U$$1799/A1 U$$1557/A2 U$$2623/A1 U$$1557/B2 VGND VGND VPWR VPWR U$$1526/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1536 U$$1536/A U$$1574/B VGND VGND VPWR VPWR U$$1536/X sky130_fd_sc_hd__xor2_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1547 U$$997/B1 U$$1557/A2 U$$864/A1 U$$1557/B2 VGND VGND VPWR VPWR U$$1548/A sky130_fd_sc_hd__a22o_1
XU$$1558 U$$1558/A U$$1558/B VGND VGND VPWR VPWR U$$1558/X sky130_fd_sc_hd__xor2_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_475 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1569 U$$3348/B1 U$$1575/A2 U$$610/B1 U$$1575/B2 VGND VGND VPWR VPWR U$$1570/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_228_ _357_/CLK _228_/D VGND VGND VPWR VPWR _228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_3 dadda_fa_2_60_3/A dadda_fa_2_60_3/B dadda_fa_2_60_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/B dadda_fa_3_60_3/B sky130_fd_sc_hd__fa_1
XFILLER_111_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater403 U$$749/A2 VGND VGND VPWR VPWR U$$739/A2 sky130_fd_sc_hd__buf_4
Xrepeater414 U$$552/X VGND VGND VPWR VPWR U$$672/A2 sky130_fd_sc_hd__buf_6
XFILLER_66_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater425 U$$521/A2 VGND VGND VPWR VPWR U$$515/A2 sky130_fd_sc_hd__buf_4
XFILLER_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_53_2 dadda_fa_2_53_2/A dadda_fa_2_53_2/B dadda_fa_2_53_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/A dadda_fa_3_53_3/A sky130_fd_sc_hd__fa_1
Xrepeater436 U$$4238/A2 VGND VGND VPWR VPWR U$$4188/A2 sky130_fd_sc_hd__buf_6
XFILLER_66_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater447 U$$4043/A2 VGND VGND VPWR VPWR U$$4011/A2 sky130_fd_sc_hd__buf_4
XFILLER_38_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4140 U$$4275/B1 U$$4164/A2 U$$4277/B1 U$$4164/B2 VGND VGND VPWR VPWR U$$4141/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater458 U$$3840/X VGND VGND VPWR VPWR U$$3970/A2 sky130_fd_sc_hd__buf_6
XU$$4151 U$$4151/A U$$4189/B VGND VGND VPWR VPWR U$$4151/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_30_1 dadda_fa_5_30_1/A dadda_fa_5_30_1/B dadda_fa_5_30_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_31_0/B dadda_fa_7_30_0/A sky130_fd_sc_hd__fa_1
Xrepeater469 U$$3703/X VGND VGND VPWR VPWR U$$3773/A2 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_46_1 U$$3158/X U$$3208/B input197/X VGND VGND VPWR VPWR dadda_fa_3_47_0/CIN
+ dadda_fa_3_46_2/CIN sky130_fd_sc_hd__fa_1
XU$$4162 U$$4162/A1 U$$4164/A2 U$$4162/B1 U$$4164/B2 VGND VGND VPWR VPWR U$$4163/A
+ sky130_fd_sc_hd__a22o_1
XU$$4173 U$$4173/A U$$4246/A VGND VGND VPWR VPWR U$$4173/X sky130_fd_sc_hd__xor2_1
XU$$4184 U$$4458/A1 U$$4226/A2 U$$4460/A1 U$$4226/B2 VGND VGND VPWR VPWR U$$4185/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_5_23_0 dadda_fa_5_23_0/A dadda_fa_5_23_0/B dadda_fa_5_23_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_24_0/A dadda_fa_6_23_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4195 U$$4195/A U$$4211/B VGND VGND VPWR VPWR U$$4195/X sky130_fd_sc_hd__xor2_1
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3450 U$$3450/A U$$3454/B VGND VGND VPWR VPWR U$$3450/X sky130_fd_sc_hd__xor2_1
XU$$3461 U$$4009/A1 U$$3479/A2 U$$3737/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3462/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_39_0 U$$1149/X U$$1282/X U$$1415/X VGND VGND VPWR VPWR dadda_fa_3_40_0/B
+ dadda_fa_3_39_2/B sky130_fd_sc_hd__fa_1
XU$$3472 U$$3472/A U$$3504/B VGND VGND VPWR VPWR U$$3472/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3483 U$$3618/B1 U$$3489/A2 U$$3483/B1 U$$3489/B2 VGND VGND VPWR VPWR U$$3484/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3494 U$$3494/A U$$3510/B VGND VGND VPWR VPWR U$$3494/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2760 U$$3719/A1 U$$2790/A2 U$$3447/A1 U$$2790/B2 VGND VGND VPWR VPWR U$$2761/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2771 U$$2771/A U$$2783/B VGND VGND VPWR VPWR U$$2771/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2782 U$$4013/B1 U$$2782/A2 U$$3878/B1 U$$2782/B2 VGND VGND VPWR VPWR U$$2783/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2793 U$$2793/A U$$2797/B VGND VGND VPWR VPWR U$$2793/X sky130_fd_sc_hd__xor2_1
XFILLER_33_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_68_2 dadda_fa_4_68_2/A dadda_fa_4_68_2/B dadda_fa_4_68_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_69_0/CIN dadda_fa_5_68_1/CIN sky130_fd_sc_hd__fa_1
Xinput206 c[54] VGND VGND VPWR VPWR input206/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput217 c[64] VGND VGND VPWR VPWR input217/X sky130_fd_sc_hd__clkbuf_1
Xinput228 c[74] VGND VGND VPWR VPWR input228/X sky130_fd_sc_hd__buf_2
XFILLER_48_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput239 c[84] VGND VGND VPWR VPWR input239/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$700 final_adder.U$$716/B final_adder.U$$700/B VGND VGND VPWR VPWR
+ final_adder.U$$780/A sky130_fd_sc_hd__and2_1
XTAP_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$711 final_adder.U$$710/B final_adder.U$$607/X final_adder.U$$591/X
+ VGND VGND VPWR VPWR final_adder.U$$711/X sky130_fd_sc_hd__a21o_1
XTAP_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_38_0 dadda_fa_7_38_0/A dadda_fa_7_38_0/B dadda_fa_7_38_0/CIN VGND VGND
+ VPWR VPWR _335_/D _206_/D sky130_fd_sc_hd__fa_2
XTAP_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$733 final_adder.U$$716/A final_adder.U$$505/X final_adder.U$$613/X
+ VGND VGND VPWR VPWR final_adder.U$$733/X sky130_fd_sc_hd__a21o_2
XTAP_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$744 final_adder.U$$776/B final_adder.U$$744/B VGND VGND VPWR VPWR
+ final_adder.U$$744/X sky130_fd_sc_hd__and2_1
XFILLER_84_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$755 final_adder.U$$754/B final_adder.U$$675/X final_adder.U$$643/X
+ VGND VGND VPWR VPWR final_adder.U$$755/X sky130_fd_sc_hd__a21o_1
XFILLER_99_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$766 final_adder.U$$798/B final_adder.U$$766/B VGND VGND VPWR VPWR
+ final_adder.U$$766/X sky130_fd_sc_hd__and2_1
XFILLER_186_1112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater970 U$$3499/A1 VGND VGND VPWR VPWR U$$896/A1 sky130_fd_sc_hd__buf_4
XU$$605 U$$605/A U$$637/B VGND VGND VPWR VPWR U$$605/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$777 final_adder.U$$776/B final_adder.U$$697/X final_adder.U$$665/X
+ VGND VGND VPWR VPWR final_adder.U$$777/X sky130_fd_sc_hd__a21o_1
Xrepeater981 U$$4456/A1 VGND VGND VPWR VPWR U$$4045/A1 sky130_fd_sc_hd__buf_8
XU$$616 U$$68/A1 U$$616/A2 U$$616/B1 U$$616/B2 VGND VGND VPWR VPWR U$$617/A sky130_fd_sc_hd__a22o_1
XFILLER_44_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$788 final_adder.U$$788/A final_adder.U$$788/B VGND VGND VPWR VPWR
+ final_adder.U$$788/X sky130_fd_sc_hd__and2_1
XFILLER_16_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$627 U$$627/A U$$673/B VGND VGND VPWR VPWR U$$627/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_1_41_0 U$$89/X U$$222/X U$$355/X VGND VGND VPWR VPWR dadda_fa_2_42_3/B dadda_fa_2_41_5/A
+ sky130_fd_sc_hd__fa_1
XFILLER_99_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_1134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater992 U$$1714/A1 VGND VGND VPWR VPWR U$$70/A1 sky130_fd_sc_hd__buf_4
XFILLER_95_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$799 final_adder.U$$798/B final_adder.U$$719/X final_adder.U$$687/X
+ VGND VGND VPWR VPWR final_adder.U$$799/X sky130_fd_sc_hd__a21o_1
XU$$638 U$$773/B1 U$$652/A2 U$$640/A1 U$$652/B2 VGND VGND VPWR VPWR U$$639/A sky130_fd_sc_hd__a22o_1
XFILLER_204_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$649 U$$649/A U$$651/B VGND VGND VPWR VPWR U$$649/X sky130_fd_sc_hd__xor2_1
XFILLER_204_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1505 input122/X VGND VGND VPWR VPWR U$$3281/A1 sky130_fd_sc_hd__buf_4
Xrepeater1516 U$$3416/A1 VGND VGND VPWR VPWR U$$2318/B1 sky130_fd_sc_hd__buf_4
XFILLER_158_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1527 input120/X VGND VGND VPWR VPWR U$$3852/B1 sky130_fd_sc_hd__buf_4
XFILLER_193_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1538 U$$3551/A1 VGND VGND VPWR VPWR U$$3414/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_158_1236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1549 U$$4369/B1 VGND VGND VPWR VPWR U$$2316/A1 sky130_fd_sc_hd__buf_4
XFILLER_125_358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_70_2 dadda_fa_3_70_2/A dadda_fa_3_70_2/B dadda_fa_3_70_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_1/A dadda_fa_4_70_2/B sky130_fd_sc_hd__fa_1
XFILLER_106_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_63_1 dadda_fa_3_63_1/A dadda_fa_3_63_1/B dadda_fa_3_63_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_0/CIN dadda_fa_4_63_2/A sky130_fd_sc_hd__fa_1
XFILLER_94_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_40_0 dadda_fa_6_40_0/A dadda_fa_6_40_0/B dadda_fa_6_40_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_41_0/B dadda_fa_7_40_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_56_0 dadda_fa_3_56_0/A dadda_fa_3_56_0/B dadda_fa_3_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_0/B dadda_fa_4_56_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_43_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2001 U$$2001/A U$$2043/B VGND VGND VPWR VPWR U$$2001/X sky130_fd_sc_hd__xor2_1
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2012 U$$2834/A1 U$$2022/A2 U$$2425/A1 U$$2022/B2 VGND VGND VPWR VPWR U$$2013/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2023 U$$2023/A U$$2037/B VGND VGND VPWR VPWR U$$2023/X sky130_fd_sc_hd__xor2_1
XFILLER_165_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2034 U$$936/B1 U$$2046/A2 U$$2445/B1 U$$2046/B2 VGND VGND VPWR VPWR U$$2035/A
+ sky130_fd_sc_hd__a22o_1
XU$$2045 U$$2045/A input22/X VGND VGND VPWR VPWR U$$2045/X sky130_fd_sc_hd__xor2_1
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1300 U$$1300/A U$$1354/B VGND VGND VPWR VPWR U$$1300/X sky130_fd_sc_hd__xor2_1
XU$$1311 U$$1448/A1 U$$1311/A2 U$$902/A1 U$$1355/B2 VGND VGND VPWR VPWR U$$1312/A
+ sky130_fd_sc_hd__a22o_1
XU$$2056 input24/X VGND VGND VPWR VPWR U$$2058/B sky130_fd_sc_hd__inv_1
XFILLER_63_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1322 U$$1322/A U$$1354/B VGND VGND VPWR VPWR U$$1322/X sky130_fd_sc_hd__xor2_1
XU$$2067 U$$2202/B1 U$$2099/A2 U$$2069/A1 U$$2099/B2 VGND VGND VPWR VPWR U$$2068/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1333 U$$2975/B1 U$$1237/X U$$2842/A1 U$$1337/B2 VGND VGND VPWR VPWR U$$1334/A
+ sky130_fd_sc_hd__a22o_1
XU$$2078 U$$2078/A U$$2094/B VGND VGND VPWR VPWR U$$2078/X sky130_fd_sc_hd__xor2_1
XU$$2089 U$$4005/B1 U$$2091/A2 U$$4009/A1 U$$2091/B2 VGND VGND VPWR VPWR U$$2090/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1344 U$$1344/A U$$1370/A VGND VGND VPWR VPWR U$$1344/X sky130_fd_sc_hd__xor2_1
XU$$1355 U$$122/A1 U$$1361/A2 U$$3547/B1 U$$1355/B2 VGND VGND VPWR VPWR U$$1356/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1366 U$$1366/A U$$1366/B VGND VGND VPWR VPWR U$$1366/X sky130_fd_sc_hd__xor2_1
XU$$1377 U$$1377/A U$$1405/B VGND VGND VPWR VPWR U$$1377/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1388 U$$1799/A1 U$$1422/A2 U$$1799/B1 U$$1422/B2 VGND VGND VPWR VPWR U$$1389/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1399 U$$1399/A U$$1399/B VGND VGND VPWR VPWR U$$1399/X sky130_fd_sc_hd__xor2_1
XFILLER_148_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_113_0 dadda_fa_7_113_0/A dadda_fa_7_113_0/B dadda_fa_7_113_0/CIN VGND
+ VGND VPWR VPWR _410_/D _281_/D sky130_fd_sc_hd__fa_1
XFILLER_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_78_1 dadda_fa_5_78_1/A dadda_fa_5_78_1/B dadda_fa_5_78_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_79_0/B dadda_fa_7_78_0/A sky130_fd_sc_hd__fa_1
XFILLER_143_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$40 _336_/Q _208_/Q VGND VGND VPWR VPWR final_adder.U$$985/B1 final_adder.U$$214/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$51 _347_/Q _219_/Q VGND VGND VPWR VPWR final_adder.U$$205/B1 final_adder.U$$204/B
+ sky130_fd_sc_hd__ha_1
XU$$3280 U$$3280/A U$$3286/B VGND VGND VPWR VPWR U$$3280/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$62 _358_/Q _230_/Q VGND VGND VPWR VPWR final_adder.U$$963/B1 final_adder.U$$192/A
+ sky130_fd_sc_hd__ha_1
XU$$3291 input44/X U$$3291/B VGND VGND VPWR VPWR U$$3291/X sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$73 _369_/Q _241_/Q VGND VGND VPWR VPWR final_adder.U$$183/B1 final_adder.U$$182/B
+ sky130_fd_sc_hd__ha_2
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$84 _380_/Q _252_/Q VGND VGND VPWR VPWR final_adder.U$$941/B1 final_adder.U$$170/A
+ sky130_fd_sc_hd__ha_1
XFILLER_94_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$95 _391_/Q _263_/Q VGND VGND VPWR VPWR final_adder.U$$161/B1 final_adder.U$$160/B
+ sky130_fd_sc_hd__ha_1
XU$$2590 U$$3547/B1 U$$2600/A2 U$$3414/A1 U$$2600/B2 VGND VGND VPWR VPWR U$$2591/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_1015 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_80_1 dadda_fa_4_80_1/A dadda_fa_4_80_1/B dadda_fa_4_80_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/B dadda_fa_5_80_1/B sky130_fd_sc_hd__fa_1
XFILLER_134_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_73_0 dadda_fa_4_73_0/A dadda_fa_4_73_0/B dadda_fa_4_73_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/A dadda_fa_5_73_1/A sky130_fd_sc_hd__fa_1
XFILLER_116_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_89_0 U$$1780/Y U$$1914/X U$$2047/X VGND VGND VPWR VPWR dadda_fa_2_90_3/CIN
+ dadda_fa_2_89_5/A sky130_fd_sc_hd__fa_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_26 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$530 final_adder.U$$538/B final_adder.U$$530/B VGND VGND VPWR VPWR
+ final_adder.U$$650/B sky130_fd_sc_hd__and2_1
XFILLER_185_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$541 final_adder.U$$540/B final_adder.U$$425/X final_adder.U$$417/X
+ VGND VGND VPWR VPWR final_adder.U$$541/X sky130_fd_sc_hd__a21o_1
XTAP_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$552 final_adder.U$$560/B final_adder.U$$552/B VGND VGND VPWR VPWR
+ final_adder.U$$672/B sky130_fd_sc_hd__and2_1
XFILLER_151_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$563 final_adder.U$$562/B final_adder.U$$447/X final_adder.U$$439/X
+ VGND VGND VPWR VPWR final_adder.U$$563/X sky130_fd_sc_hd__a21o_1
XTAP_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$402 U$$676/A1 U$$278/X U$$676/B1 U$$279/X VGND VGND VPWR VPWR U$$403/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$574 final_adder.U$$582/B final_adder.U$$574/B VGND VGND VPWR VPWR
+ final_adder.U$$694/B sky130_fd_sc_hd__and2_1
XTAP_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$413 U$$536/B VGND VGND VPWR VPWR U$$413/Y sky130_fd_sc_hd__inv_1
XFILLER_56_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$585 final_adder.U$$584/B final_adder.U$$469/X final_adder.U$$461/X
+ VGND VGND VPWR VPWR final_adder.U$$585/X sky130_fd_sc_hd__a21o_1
XU$$424 U$$424/A U$$436/B VGND VGND VPWR VPWR U$$424/X sky130_fd_sc_hd__xor2_1
XTAP_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$596 final_adder.U$$604/B final_adder.U$$596/B VGND VGND VPWR VPWR
+ final_adder.U$$716/B sky130_fd_sc_hd__and2_1
XU$$435 U$$24/A1 U$$515/A2 U$$26/A1 U$$515/B2 VGND VGND VPWR VPWR U$$436/A sky130_fd_sc_hd__a22o_1
XTAP_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_76 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$446 U$$446/A U$$516/B VGND VGND VPWR VPWR U$$446/X sky130_fd_sc_hd__xor2_1
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$457 U$$594/A1 U$$491/A2 U$$594/B1 U$$491/B2 VGND VGND VPWR VPWR U$$458/A sky130_fd_sc_hd__a22o_1
XFILLER_72_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$468 U$$468/A U$$484/B VGND VGND VPWR VPWR U$$468/X sky130_fd_sc_hd__xor2_1
XU$$479 U$$68/A1 U$$483/A2 U$$616/B1 U$$483/B2 VGND VGND VPWR VPWR U$$480/A sky130_fd_sc_hd__a22o_1
XFILLER_71_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_88_0 dadda_fa_6_88_0/A dadda_fa_6_88_0/B dadda_fa_6_88_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_89_0/B dadda_fa_7_88_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1302 input47/X VGND VGND VPWR VPWR U$$3510/B sky130_fd_sc_hd__buf_6
XFILLER_154_954 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1313 U$$3244/B VGND VGND VPWR VPWR U$$3208/B sky130_fd_sc_hd__buf_8
XFILLER_126_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1324 U$$3151/A VGND VGND VPWR VPWR U$$3109/B sky130_fd_sc_hd__buf_6
Xdadda_ha_0_78_0 dadda_ha_0_78_0/A U$$1094/X VGND VGND VPWR VPWR dadda_fa_2_79_0/A
+ dadda_fa_2_78_0/A sky130_fd_sc_hd__ha_1
Xrepeater1335 input38/X VGND VGND VPWR VPWR U$$2978/B sky130_fd_sc_hd__buf_6
XFILLER_126_667 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1346 U$$2845/B VGND VGND VPWR VPWR U$$2876/A sky130_fd_sc_hd__buf_6
XFILLER_4_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1357 U$$274/A VGND VGND VPWR VPWR U$$272/B sky130_fd_sc_hd__clkbuf_8
XFILLER_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1368 U$$2603/A VGND VGND VPWR VPWR U$$2602/A sky130_fd_sc_hd__buf_6
XFILLER_119_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1379 U$$808/B VGND VGND VPWR VPWR U$$821/A sky130_fd_sc_hd__buf_8
XFILLER_84_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4465_1809 VGND VGND VPWR VPWR U$$4465_1809/HI U$$4465/B sky130_fd_sc_hd__conb_1
XFILLER_48_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_1012 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1056 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$980 U$$980/A U$$980/B VGND VGND VPWR VPWR U$$980/X sky130_fd_sc_hd__xor2_1
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$991 U$$991/A1 U$$993/A2 U$$993/A1 U$$993/B2 VGND VGND VPWR VPWR U$$992/A sky130_fd_sc_hd__a22o_1
XU$$1130 U$$2363/A1 U$$1136/A2 U$$995/A1 U$$1136/B2 VGND VGND VPWR VPWR U$$1131/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1141 U$$1141/A U$$1175/B VGND VGND VPWR VPWR U$$1141/X sky130_fd_sc_hd__xor2_1
XU$$1152 U$$328/B1 U$$1162/A2 U$$58/A1 U$$1162/B2 VGND VGND VPWR VPWR U$$1153/A sky130_fd_sc_hd__a22o_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1163 U$$1163/A U$$1195/B VGND VGND VPWR VPWR U$$1163/X sky130_fd_sc_hd__xor2_1
XFILLER_206_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1174 U$$1448/A1 U$$1174/A2 U$$902/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1175/A
+ sky130_fd_sc_hd__a22o_1
XU$$1185 U$$1185/A U$$1223/B VGND VGND VPWR VPWR U$$1185/X sky130_fd_sc_hd__xor2_1
XFILLER_203_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1196 U$$98/B1 U$$1204/A2 U$$924/A1 U$$1204/B2 VGND VGND VPWR VPWR U$$1197/A sky130_fd_sc_hd__a22o_1
XFILLER_52_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_90_0 dadda_fa_5_90_0/A dadda_fa_5_90_0/B dadda_fa_5_90_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_91_0/A dadda_fa_6_90_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_75_6 U$$4014/X U$$4147/X U$$4280/X VGND VGND VPWR VPWR dadda_fa_2_76_2/B
+ dadda_fa_2_75_5/B sky130_fd_sc_hd__fa_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_68_5 input221/X dadda_fa_1_68_5/B dadda_fa_1_68_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_69_2/A dadda_fa_2_68_5/A sky130_fd_sc_hd__fa_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 _384_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_119 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_120_0 dadda_fa_6_120_0/A dadda_fa_6_120_0/B dadda_fa_6_120_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_121_0/B dadda_fa_7_120_0/CIN sky130_fd_sc_hd__fa_1
XTAP_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_63_4 U$$1729/X U$$1862/X U$$1995/X VGND VGND VPWR VPWR dadda_fa_1_64_6/CIN
+ dadda_fa_1_63_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_40_3 dadda_fa_3_40_3/A dadda_fa_3_40_3/B dadda_fa_3_40_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_41_1/B dadda_fa_4_40_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$360 final_adder.U$$362/B final_adder.U$$360/B VGND VGND VPWR VPWR
+ final_adder.U$$486/B sky130_fd_sc_hd__and2_1
XTAP_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$371 final_adder.U$$370/B final_adder.U$$245/X final_adder.U$$243/X
+ VGND VGND VPWR VPWR final_adder.U$$371/X sky130_fd_sc_hd__a21o_1
XTAP_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$210 U$$210/A U$$212/B VGND VGND VPWR VPWR U$$210/X sky130_fd_sc_hd__xor2_1
XTAP_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$221 U$$630/B1 U$$263/A2 U$$86/A1 U$$231/B2 VGND VGND VPWR VPWR U$$222/A sky130_fd_sc_hd__a22o_1
XFILLER_57_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_33_2 dadda_fa_3_33_2/A dadda_fa_3_33_2/B dadda_fa_3_33_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_1/A dadda_fa_4_33_2/B sky130_fd_sc_hd__fa_1
XTAP_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$393 final_adder.U$$392/B final_adder.U$$271/X final_adder.U$$267/X
+ VGND VGND VPWR VPWR final_adder.U$$393/X sky130_fd_sc_hd__a21o_1
XTAP_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$232 U$$232/A U$$264/B VGND VGND VPWR VPWR U$$232/X sky130_fd_sc_hd__xor2_1
XFILLER_40_1188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$243 U$$654/A1 U$$243/A2 U$$654/B1 U$$243/B2 VGND VGND VPWR VPWR U$$244/A sky130_fd_sc_hd__a22o_1
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$254 U$$254/A U$$260/B VGND VGND VPWR VPWR U$$254/X sky130_fd_sc_hd__xor2_1
XTAP_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$265 U$$676/A1 U$$141/X U$$676/B1 U$$142/X VGND VGND VPWR VPWR U$$266/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_26_1 U$$1522/X U$$1655/X U$$1788/X VGND VGND VPWR VPWR dadda_fa_4_27_0/CIN
+ dadda_fa_4_26_2/A sky130_fd_sc_hd__fa_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$276 U$$411/A VGND VGND VPWR VPWR U$$276/Y sky130_fd_sc_hd__inv_1
XU$$287 U$$287/A U$$317/B VGND VGND VPWR VPWR U$$287/X sky130_fd_sc_hd__xor2_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$298 U$$24/A1 U$$302/A2 U$$26/A1 U$$302/B2 VGND VGND VPWR VPWR U$$299/A sky130_fd_sc_hd__a22o_1
XFILLER_72_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_19_0 U$$45/X U$$178/X U$$311/X VGND VGND VPWR VPWR dadda_fa_4_20_0/CIN
+ dadda_fa_4_19_2/A sky130_fd_sc_hd__fa_1
XFILLER_44_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4 U$$2/Y U$$1/A U$$4/A3 U$$3/X U$$0/Y VGND VGND VPWR VPWR U$$4/X sky130_fd_sc_hd__a32o_1
XFILLER_51_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1019 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1110 U$$44/B1 VGND VGND VPWR VPWR U$$46/A1 sky130_fd_sc_hd__buf_4
Xrepeater1121 input74/X VGND VGND VPWR VPWR U$$4428/A1 sky130_fd_sc_hd__buf_4
Xoutput307 output307/A VGND VGND VPWR VPWR o[2] sky130_fd_sc_hd__buf_2
XFILLER_160_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput318 output318/A VGND VGND VPWR VPWR o[3] sky130_fd_sc_hd__buf_2
Xrepeater1132 input72/X VGND VGND VPWR VPWR U$$38/B1 sky130_fd_sc_hd__clkbuf_8
Xoutput329 output329/A VGND VGND VPWR VPWR o[4] sky130_fd_sc_hd__buf_2
XFILLER_154_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1143 U$$3737/A1 VGND VGND VPWR VPWR U$$860/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1154 U$$1076/B VGND VGND VPWR VPWR U$$994/B sky130_fd_sc_hd__buf_6
XFILLER_114_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_85_5 dadda_fa_2_85_5/A dadda_fa_2_85_5/B dadda_fa_2_85_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_86_2/A dadda_fa_4_85_0/A sky130_fd_sc_hd__fa_2
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1165 U$$2363/A1 VGND VGND VPWR VPWR U$$993/A1 sky130_fd_sc_hd__buf_4
XFILLER_141_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1176 U$$4005/A1 VGND VGND VPWR VPWR U$$4277/B1 sky130_fd_sc_hd__buf_6
Xrepeater1187 input67/X VGND VGND VPWR VPWR U$$4275/B1 sky130_fd_sc_hd__buf_6
Xrepeater1198 U$$1515/A1 VGND VGND VPWR VPWR U$$967/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_141_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_78_4 dadda_fa_2_78_4/A dadda_fa_2_78_4/B dadda_fa_2_78_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_1/CIN dadda_fa_3_78_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_101_3 U$$3800/X U$$3933/X U$$4066/X VGND VGND VPWR VPWR dadda_fa_3_102_2/CIN
+ dadda_fa_4_101_0/A sky130_fd_sc_hd__fa_1
XFILLER_91_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_115_1 dadda_fa_5_115_1/A dadda_fa_5_115_1/B dadda_fa_5_115_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_116_0/B dadda_fa_7_115_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_108_0 dadda_fa_5_108_0/A dadda_fa_5_108_0/B dadda_fa_5_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_109_0/A dadda_fa_6_108_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_80_4 U$$2694/X U$$2827/X U$$2960/X VGND VGND VPWR VPWR dadda_fa_2_81_2/A
+ dadda_fa_2_80_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_73_3 U$$3079/X U$$3212/X U$$3345/X VGND VGND VPWR VPWR dadda_fa_2_74_1/B
+ dadda_fa_2_73_4/B sky130_fd_sc_hd__fa_1
XFILLER_141_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_50_2 dadda_fa_4_50_2/A dadda_fa_4_50_2/B dadda_fa_4_50_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_51_0/CIN dadda_fa_5_50_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4487_1820 VGND VGND VPWR VPWR U$$4487_1820/HI U$$4487/B sky130_fd_sc_hd__conb_1
Xdadda_fa_1_66_2 U$$3331/X U$$3464/X U$$3597/X VGND VGND VPWR VPWR dadda_fa_2_67_1/A
+ dadda_fa_2_66_4/A sky130_fd_sc_hd__fa_1
XFILLER_59_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_43_1 dadda_fa_4_43_1/A dadda_fa_4_43_1/B dadda_fa_4_43_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/B dadda_fa_5_43_1/B sky130_fd_sc_hd__fa_1
XFILLER_111_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_59_1 U$$1987/X U$$2120/X U$$2253/X VGND VGND VPWR VPWR dadda_fa_2_60_0/CIN
+ dadda_fa_2_59_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_7_20_0 dadda_fa_7_20_0/A dadda_fa_7_20_0/B dadda_fa_7_20_0/CIN VGND VGND
+ VPWR VPWR _317_/D _188_/D sky130_fd_sc_hd__fa_1
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_36_0 dadda_fa_4_36_0/A dadda_fa_4_36_0/B dadda_fa_4_36_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/A dadda_fa_5_36_1/A sky130_fd_sc_hd__fa_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_330_ _337_/CLK _330_/D VGND VGND VPWR VPWR _330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _381_/CLK _261_/D VGND VGND VPWR VPWR _261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_192_ _329_/CLK _192_/D VGND VGND VPWR VPWR _192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_88_3 dadda_fa_3_88_3/A dadda_fa_3_88_3/B dadda_fa_3_88_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_89_1/B dadda_fa_4_88_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_543 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4503 U$$4503/A U$$4503/B VGND VGND VPWR VPWR U$$4503/X sky130_fd_sc_hd__xor2_1
XU$$4514 U$$4514/A1 U$$4388/X U$$4516/A1 U$$4389/X VGND VGND VPWR VPWR U$$4515/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_0_61_1 U$$528/X U$$661/X U$$794/X VGND VGND VPWR VPWR dadda_fa_1_62_6/A
+ dadda_fa_1_61_8/A sky130_fd_sc_hd__fa_1
XTAP_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3802 U$$3802/A U$$3814/B VGND VGND VPWR VPWR U$$3802/X sky130_fd_sc_hd__xor2_1
XU$$17 U$$17/A U$$9/B VGND VGND VPWR VPWR U$$17/X sky130_fd_sc_hd__xor2_1
XTAP_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$28 U$$28/A1 U$$50/A2 U$$30/A1 U$$50/B2 VGND VGND VPWR VPWR U$$29/A sky130_fd_sc_hd__a22o_1
XU$$3813 U$$3813/A1 U$$3813/A2 U$$388/B1 U$$3813/B2 VGND VGND VPWR VPWR U$$3814/A
+ sky130_fd_sc_hd__a22o_1
XU$$3824 U$$3824/A U$$3826/B VGND VGND VPWR VPWR U$$3824/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_54_0 U$$115/X U$$248/X U$$381/X VGND VGND VPWR VPWR dadda_fa_1_55_8/A
+ dadda_fa_1_54_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$39 U$$39/A U$$43/B VGND VGND VPWR VPWR U$$39/X sky130_fd_sc_hd__xor2_1
XU$$3835 U$$3836/A VGND VGND VPWR VPWR U$$3835/Y sky130_fd_sc_hd__inv_1
XTAP_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3846 input76/X U$$3878/A2 U$$3846/B1 U$$3878/B2 VGND VGND VPWR VPWR U$$3847/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$190 final_adder.U$$190/A final_adder.U$$190/B VGND VGND VPWR VPWR
+ final_adder.U$$318/B sky130_fd_sc_hd__and2_1
XTAP_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3857 U$$3857/A U$$3875/B VGND VGND VPWR VPWR U$$3857/X sky130_fd_sc_hd__xor2_1
XFILLER_79_1151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3868 U$$4277/B1 U$$3902/A2 U$$4418/A1 U$$3902/B2 VGND VGND VPWR VPWR U$$3869/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3879 U$$3879/A U$$3879/B VGND VGND VPWR VPWR U$$3879/X sky130_fd_sc_hd__xor2_1
XTAP_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 _336_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_202_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1010 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_90_3 U$$4443/X input246/X dadda_fa_2_90_3/CIN VGND VGND VPWR VPWR dadda_fa_3_91_1/B
+ dadda_fa_3_90_3/B sky130_fd_sc_hd__fa_1
XFILLER_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_83_2 dadda_fa_2_83_2/A dadda_fa_2_83_2/B dadda_fa_2_83_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/A dadda_fa_3_83_3/A sky130_fd_sc_hd__fa_1
XFILLER_82_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1019 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_60_1 dadda_fa_5_60_1/A dadda_fa_5_60_1/B dadda_fa_5_60_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_61_0/B dadda_fa_7_60_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_76_1 dadda_fa_2_76_1/A dadda_fa_2_76_1/B dadda_fa_2_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_0/CIN dadda_fa_3_76_2/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_5_53_0 dadda_fa_5_53_0/A dadda_fa_5_53_0/B dadda_fa_5_53_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_54_0/A dadda_fa_6_53_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_830 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_69_0 dadda_fa_2_69_0/A dadda_fa_2_69_0/B dadda_fa_2_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_0/B dadda_fa_3_69_2/B sky130_fd_sc_hd__fa_1
XFILLER_110_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_885 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_52_8 U$$3569/X U$$3609/B input204/X VGND VGND VPWR VPWR dadda_fa_2_53_3/A
+ dadda_fa_3_52_0/A sky130_fd_sc_hd__fa_2
XFILLER_3_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_410 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_98_2 dadda_fa_4_98_2/A dadda_fa_4_98_2/B dadda_fa_4_98_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_99_0/CIN dadda_fa_5_98_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_194_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_68_0 dadda_fa_7_68_0/A dadda_fa_7_68_0/B dadda_fa_7_68_0/CIN VGND VGND
+ VPWR VPWR _365_/D _236_/D sky130_fd_sc_hd__fa_1
XFILLER_65_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_71_0 U$$2144/X U$$2277/X U$$2410/X VGND VGND VPWR VPWR dadda_fa_2_72_0/B
+ dadda_fa_2_71_3/B sky130_fd_sc_hd__fa_1
XFILLER_114_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3109 U$$3109/A U$$3109/B VGND VGND VPWR VPWR U$$3109/X sky130_fd_sc_hd__xor2_1
XFILLER_100_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2408 U$$2408/A U$$2446/B VGND VGND VPWR VPWR U$$2408/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1029 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2419 U$$3787/B1 U$$2459/A2 U$$914/A1 U$$2459/B2 VGND VGND VPWR VPWR U$$2420/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1707 U$$1707/A U$$1707/B VGND VGND VPWR VPWR U$$1707/X sky130_fd_sc_hd__xor2_1
XFILLER_28_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1718 U$$483/B1 U$$1750/A2 U$$2951/B1 U$$1750/B2 VGND VGND VPWR VPWR U$$1719/A
+ sky130_fd_sc_hd__a22o_1
XU$$1729 U$$1729/A U$$1739/B VGND VGND VPWR VPWR U$$1729/X sky130_fd_sc_hd__xor2_1
XFILLER_42_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_313_ _314_/CLK _313_/D VGND VGND VPWR VPWR _313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1002 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_244_ _373_/CLK _244_/D VGND VGND VPWR VPWR _244_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_167_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput17 a[24] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput28 a[34] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 a[44] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_1
X_175_ _327_/CLK _175_/D VGND VGND VPWR VPWR _175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_93_1 dadda_fa_3_93_1/A dadda_fa_3_93_1/B dadda_fa_3_93_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_0/CIN dadda_fa_4_93_2/A sky130_fd_sc_hd__fa_1
XFILLER_182_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_70_0 dadda_fa_6_70_0/A dadda_fa_6_70_0/B dadda_fa_6_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_71_0/B dadda_fa_7_70_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_86_0 dadda_fa_3_86_0/A dadda_fa_3_86_0/B dadda_fa_3_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_0/B dadda_fa_4_86_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater607 U$$1511/X VGND VGND VPWR VPWR U$$1637/A2 sky130_fd_sc_hd__buf_6
XU$$4300 U$$4300/A U$$4384/A VGND VGND VPWR VPWR U$$4300/X sky130_fd_sc_hd__xor2_1
Xrepeater618 U$$1422/A2 VGND VGND VPWR VPWR U$$1404/A2 sky130_fd_sc_hd__clkbuf_4
Xrepeater629 U$$1237/X VGND VGND VPWR VPWR U$$1337/A2 sky130_fd_sc_hd__buf_4
XFILLER_77_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4311 U$$4311/A1 U$$4369/A2 U$$4311/B1 U$$4369/B2 VGND VGND VPWR VPWR U$$4312/A
+ sky130_fd_sc_hd__a22o_1
XU$$4322 U$$4322/A U$$4330/B VGND VGND VPWR VPWR U$$4322/X sky130_fd_sc_hd__xor2_1
XU$$4333 U$$4333/A1 U$$4349/A2 U$$4333/B1 U$$4349/B2 VGND VGND VPWR VPWR U$$4334/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4344 U$$4344/A U$$4354/B VGND VGND VPWR VPWR U$$4344/X sky130_fd_sc_hd__xor2_1
XFILLER_133_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4355 U$$4492/A1 U$$4361/A2 U$$4494/A1 U$$4361/B2 VGND VGND VPWR VPWR U$$4356/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3610 U$$4293/B1 U$$3644/A2 U$$3884/B1 U$$3644/B2 VGND VGND VPWR VPWR U$$3611/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_115_0 U$$3961/X U$$4094/X U$$4227/X VGND VGND VPWR VPWR dadda_fa_5_116_0/A
+ dadda_fa_5_115_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_48_5 dadda_fa_2_48_5/A dadda_fa_2_48_5/B dadda_fa_2_48_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_49_2/A dadda_fa_4_48_0/A sky130_fd_sc_hd__fa_2
XU$$3621 U$$3621/A U$$3623/B VGND VGND VPWR VPWR U$$3621/X sky130_fd_sc_hd__xor2_1
XU$$4366 U$$4366/A U$$4366/B VGND VGND VPWR VPWR U$$4366/X sky130_fd_sc_hd__xor2_1
XFILLER_19_963 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3632 U$$4043/A1 U$$3636/A2 U$$4043/B1 U$$3636/B2 VGND VGND VPWR VPWR U$$3633/A
+ sky130_fd_sc_hd__a22o_1
XU$$4377 U$$4514/A1 U$$4251/X U$$4516/A1 U$$4252/X VGND VGND VPWR VPWR U$$4378/A sky130_fd_sc_hd__a22o_1
XU$$4388 U$$4386/Y U$$4388/A2 U$$4384/A U$$4387/X U$$4384/Y VGND VGND VPWR VPWR U$$4388/X
+ sky130_fd_sc_hd__a32o_1
XU$$3643 U$$3643/A U$$3643/B VGND VGND VPWR VPWR U$$3643/X sky130_fd_sc_hd__xor2_1
XFILLER_65_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3654 U$$914/A1 U$$3660/A2 U$$914/B1 U$$3660/B2 VGND VGND VPWR VPWR U$$3655/A sky130_fd_sc_hd__a22o_1
XU$$4399 U$$4399/A U$$4399/B VGND VGND VPWR VPWR U$$4399/X sky130_fd_sc_hd__xor2_1
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3665 U$$3665/A U$$3665/B VGND VGND VPWR VPWR U$$3665/X sky130_fd_sc_hd__xor2_1
XU$$2920 U$$2920/A U$$2920/B VGND VGND VPWR VPWR U$$2920/X sky130_fd_sc_hd__xor2_1
XU$$2931 U$$4438/A1 U$$2977/A2 U$$4440/A1 U$$2979/B2 VGND VGND VPWR VPWR U$$2932/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3676 U$$3813/A1 U$$3680/A2 U$$116/A1 U$$3680/B2 VGND VGND VPWR VPWR U$$3677/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3687 U$$3687/A U$$3698/A VGND VGND VPWR VPWR U$$3687/X sky130_fd_sc_hd__xor2_1
XFILLER_46_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2942 U$$2942/A U$$2950/B VGND VGND VPWR VPWR U$$2942/X sky130_fd_sc_hd__xor2_1
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3698 U$$3698/A VGND VGND VPWR VPWR U$$3698/Y sky130_fd_sc_hd__inv_1
XU$$2953 U$$3499/B1 U$$2995/A2 U$$2955/A1 U$$2995/B2 VGND VGND VPWR VPWR U$$2954/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2964 U$$2964/A input38/X VGND VGND VPWR VPWR U$$2964/X sky130_fd_sc_hd__xor2_1
XU$$2975 U$$2975/A1 U$$2977/A2 U$$2975/B1 U$$2979/B2 VGND VGND VPWR VPWR U$$2976/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2986 U$$2986/A U$$3008/B VGND VGND VPWR VPWR U$$2986/X sky130_fd_sc_hd__xor2_1
XFILLER_34_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2997 U$$3545/A1 U$$3011/A2 U$$3684/A1 U$$3011/B2 VGND VGND VPWR VPWR U$$2998/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_927 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$915 final_adder.U$$144/A final_adder.U$$853/X final_adder.U$$915/B1
+ VGND VGND VPWR VPWR final_adder.U$$915/X sky130_fd_sc_hd__a21o_1
XFILLER_151_1264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$937 final_adder.U$$166/A final_adder.U$$875/X final_adder.U$$937/B1
+ VGND VGND VPWR VPWR final_adder.U$$937/X sky130_fd_sc_hd__a21o_1
XFILLER_96_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_50_5 U$$2102/X U$$2235/X U$$2368/X VGND VGND VPWR VPWR dadda_fa_2_51_2/A
+ dadda_fa_2_50_5/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$959 final_adder.U$$188/A final_adder.U$$897/X final_adder.U$$959/B1
+ VGND VGND VPWR VPWR final_adder.U$$959/X sky130_fd_sc_hd__a21o_1
XFILLER_83_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$809 U$$944/B1 U$$689/X U$$811/A1 U$$690/X VGND VGND VPWR VPWR U$$810/A sky130_fd_sc_hd__a22o_1
XFILLER_95_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1035 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_693 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2205 U$$2205/A U$$2253/B VGND VGND VPWR VPWR U$$2205/X sky130_fd_sc_hd__xor2_1
XFILLER_207_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2216 U$$2625/B1 U$$2272/A2 U$$2492/A1 U$$2272/B2 VGND VGND VPWR VPWR U$$2217/A
+ sky130_fd_sc_hd__a22o_1
XU$$2227 U$$2227/A U$$2227/B VGND VGND VPWR VPWR U$$2227/X sky130_fd_sc_hd__xor2_1
XFILLER_90_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2238 U$$44/B1 U$$2284/A2 U$$3882/B1 U$$2284/B2 VGND VGND VPWR VPWR U$$2239/A sky130_fd_sc_hd__a22o_1
XFILLER_76_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2249 U$$2249/A U$$2285/B VGND VGND VPWR VPWR U$$2249/X sky130_fd_sc_hd__xor2_1
XU$$1504 U$$1504/A1 U$$1504/A2 U$$1504/B1 U$$1504/B2 VGND VGND VPWR VPWR U$$1505/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1515 U$$1515/A1 U$$1575/A2 U$$2202/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1516/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1526 U$$1526/A U$$1558/B VGND VGND VPWR VPWR U$$1526/X sky130_fd_sc_hd__xor2_1
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1537 U$$850/B1 U$$1575/A2 U$$854/A1 U$$1575/B2 VGND VGND VPWR VPWR U$$1538/A sky130_fd_sc_hd__a22o_1
XFILLER_188_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1548 U$$1548/A U$$1558/B VGND VGND VPWR VPWR U$$1548/X sky130_fd_sc_hd__xor2_1
XFILLER_187_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1559 U$$461/B1 U$$1591/A2 U$$328/A1 U$$1591/B2 VGND VGND VPWR VPWR U$$1560/A sky130_fd_sc_hd__a22o_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_227_ _227_/CLK _227_/D VGND VGND VPWR VPWR _227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_1174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_2_60_4 dadda_fa_2_60_4/A dadda_fa_2_60_4/B dadda_fa_2_60_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_1/CIN dadda_fa_3_60_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_97_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater404 U$$759/A2 VGND VGND VPWR VPWR U$$749/A2 sky130_fd_sc_hd__buf_6
Xrepeater415 U$$4297/A2 VGND VGND VPWR VPWR U$$4275/A2 sky130_fd_sc_hd__buf_6
Xrepeater426 U$$527/A2 VGND VGND VPWR VPWR U$$521/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_53_3 dadda_fa_2_53_3/A dadda_fa_2_53_3/B dadda_fa_2_53_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/B dadda_fa_3_53_3/B sky130_fd_sc_hd__fa_1
Xrepeater437 U$$4240/A2 VGND VGND VPWR VPWR U$$4238/A2 sky130_fd_sc_hd__buf_6
Xrepeater448 U$$4043/A2 VGND VGND VPWR VPWR U$$4035/A2 sky130_fd_sc_hd__buf_6
XFILLER_211_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater459 U$$3926/A2 VGND VGND VPWR VPWR U$$3946/A2 sky130_fd_sc_hd__buf_6
XU$$4130 U$$4402/B1 U$$4164/A2 U$$4406/A1 U$$4164/B2 VGND VGND VPWR VPWR U$$4131/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4141 U$$4141/A U$$4165/B VGND VGND VPWR VPWR U$$4141/X sky130_fd_sc_hd__xor2_1
XFILLER_38_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4152 input73/X U$$4188/A2 input74/X U$$4188/B2 VGND VGND VPWR VPWR U$$4153/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_46_2 dadda_fa_2_46_2/A dadda_fa_2_46_2/B dadda_fa_2_46_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/A dadda_fa_3_46_3/A sky130_fd_sc_hd__fa_1
XFILLER_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4163 U$$4163/A U$$4165/B VGND VGND VPWR VPWR U$$4163/X sky130_fd_sc_hd__xor2_1
XU$$4174 U$$4309/B1 U$$4176/A2 U$$4176/A1 U$$4176/B2 VGND VGND VPWR VPWR U$$4175/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3440 U$$3440/A U$$3528/B VGND VGND VPWR VPWR U$$3440/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4185 U$$4185/A U$$4227/B VGND VGND VPWR VPWR U$$4185/X sky130_fd_sc_hd__xor2_1
XFILLER_19_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_23_1 dadda_fa_5_23_1/A dadda_fa_5_23_1/B dadda_fa_5_23_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_24_0/B dadda_fa_7_23_0/A sky130_fd_sc_hd__fa_1
XU$$4196 U$$4333/A1 U$$4210/A2 U$$4333/B1 U$$4210/B2 VGND VGND VPWR VPWR U$$4197/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_39_1 U$$1548/X U$$1681/X U$$1814/X VGND VGND VPWR VPWR dadda_fa_3_40_0/CIN
+ dadda_fa_3_39_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_53_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3451 U$$3451/A1 U$$3453/A2 U$$4410/B1 U$$3453/B2 VGND VGND VPWR VPWR U$$3452/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3462 U$$3462/A U$$3480/B VGND VGND VPWR VPWR U$$3462/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3473 U$$3473/A1 U$$3479/A2 U$$3884/B1 U$$3479/B2 VGND VGND VPWR VPWR U$$3474/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3484 U$$3484/A U$$3490/B VGND VGND VPWR VPWR U$$3484/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_16_0 dadda_fa_5_16_0/A dadda_fa_5_16_0/B dadda_fa_5_16_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_17_0/A dadda_fa_6_16_0/CIN sky130_fd_sc_hd__fa_1
XU$$2750 U$$3159/B1 U$$2796/A2 U$$3026/A1 U$$2796/B2 VGND VGND VPWR VPWR U$$2751/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3495 U$$4043/A1 U$$3429/X U$$4045/A1 U$$3430/X VGND VGND VPWR VPWR U$$3496/A sky130_fd_sc_hd__a22o_1
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2761 U$$2761/A U$$2797/B VGND VGND VPWR VPWR U$$2761/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2772 U$$32/A1 U$$2782/A2 U$$32/B1 U$$2782/B2 VGND VGND VPWR VPWR U$$2773/A sky130_fd_sc_hd__a22o_1
XU$$2783 U$$2783/A U$$2783/B VGND VGND VPWR VPWR U$$2783/X sky130_fd_sc_hd__xor2_1
XFILLER_209_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2794 U$$4162/B1 U$$2796/A2 U$$3344/A1 U$$2796/B2 VGND VGND VPWR VPWR U$$2795/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput207 c[55] VGND VGND VPWR VPWR input207/X sky130_fd_sc_hd__clkbuf_4
Xinput218 c[65] VGND VGND VPWR VPWR input218/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput229 c[75] VGND VGND VPWR VPWR input229/X sky130_fd_sc_hd__buf_2
XFILLER_124_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$701 final_adder.U$$700/B final_adder.U$$597/X final_adder.U$$581/X
+ VGND VGND VPWR VPWR final_adder.U$$701/X sky130_fd_sc_hd__a21o_1
XFILLER_64_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$712 final_adder.U$$712/A final_adder.U$$712/B VGND VGND VPWR VPWR
+ final_adder.U$$792/A sky130_fd_sc_hd__and2_1
XTAP_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$723 final_adder.U$$706/A final_adder.U$$619/X final_adder.U$$603/X
+ VGND VGND VPWR VPWR final_adder.U$$723/X sky130_fd_sc_hd__a21o_2
XTAP_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$745 final_adder.U$$744/B final_adder.U$$665/X final_adder.U$$633/X
+ VGND VGND VPWR VPWR final_adder.U$$745/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$756 final_adder.U$$788/B final_adder.U$$756/B VGND VGND VPWR VPWR
+ final_adder.U$$756/X sky130_fd_sc_hd__and2_1
XFILLER_151_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater960 U$$2951/B1 VGND VGND VPWR VPWR U$$1446/A1 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$767 final_adder.U$$766/B final_adder.U$$687/X final_adder.U$$655/X
+ VGND VGND VPWR VPWR final_adder.U$$767/X sky130_fd_sc_hd__a21o_1
XFILLER_72_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater971 U$$3088/A1 VGND VGND VPWR VPWR U$$3499/A1 sky130_fd_sc_hd__buf_6
XU$$606 U$$878/B1 U$$606/A2 U$$745/A1 U$$606/B2 VGND VGND VPWR VPWR U$$607/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$778 final_adder.U$$778/A final_adder.U$$778/B VGND VGND VPWR VPWR
+ final_adder.U$$778/X sky130_fd_sc_hd__and2_1
XFILLER_186_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater982 input90/X VGND VGND VPWR VPWR U$$4456/A1 sky130_fd_sc_hd__clkbuf_8
XU$$617 U$$617/A U$$617/B VGND VGND VPWR VPWR U$$617/X sky130_fd_sc_hd__xor2_1
XFILLER_56_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$789 final_adder.U$$788/B final_adder.U$$709/X final_adder.U$$677/X
+ VGND VGND VPWR VPWR final_adder.U$$789/X sky130_fd_sc_hd__a21o_1
Xrepeater993 U$$1714/A1 VGND VGND VPWR VPWR U$$616/B1 sky130_fd_sc_hd__buf_6
XU$$628 U$$763/B1 U$$672/A2 U$$630/A1 U$$668/B2 VGND VGND VPWR VPWR U$$629/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_41_1 U$$488/X U$$621/X U$$754/X VGND VGND VPWR VPWR dadda_fa_2_42_3/CIN
+ dadda_fa_2_41_5/B sky130_fd_sc_hd__fa_1
XFILLER_112_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$639 U$$639/A U$$651/B VGND VGND VPWR VPWR U$$639/X sky130_fd_sc_hd__xor2_1
XFILLER_186_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_777 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1506 U$$950/B1 VGND VGND VPWR VPWR U$$676/B1 sky130_fd_sc_hd__buf_4
XFILLER_123_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1517 U$$3416/A1 VGND VGND VPWR VPWR U$$3414/B1 sky130_fd_sc_hd__buf_6
XFILLER_153_635 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1528 input120/X VGND VGND VPWR VPWR U$$3578/B1 sky130_fd_sc_hd__buf_6
XFILLER_119_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1539 U$$811/A1 VGND VGND VPWR VPWR U$$674/A1 sky130_fd_sc_hd__buf_4
XFILLER_193_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_808 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_70_3 dadda_fa_3_70_3/A dadda_fa_3_70_3/B dadda_fa_3_70_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_71_1/B dadda_fa_4_70_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_63_2 dadda_fa_3_63_2/A dadda_fa_3_63_2/B dadda_fa_3_63_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_1/A dadda_fa_4_63_2/B sky130_fd_sc_hd__fa_1
Xdadda_fa_3_56_1 dadda_fa_3_56_1/A dadda_fa_3_56_1/B dadda_fa_3_56_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_0/CIN dadda_fa_4_56_2/A sky130_fd_sc_hd__fa_1
XFILLER_130_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_33_0 dadda_fa_6_33_0/A dadda_fa_6_33_0/B dadda_fa_6_33_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_34_0/B dadda_fa_7_33_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_49_0 dadda_fa_3_49_0/A dadda_fa_3_49_0/B dadda_fa_3_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_0/B dadda_fa_4_49_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_207_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2002 U$$3235/A1 U$$2022/A2 U$$2415/A1 U$$2022/B2 VGND VGND VPWR VPWR U$$2003/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2013 U$$2013/A U$$2037/B VGND VGND VPWR VPWR U$$2013/X sky130_fd_sc_hd__xor2_1
XU$$2024 U$$928/A1 U$$2052/A2 U$$930/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2025/A sky130_fd_sc_hd__a22o_1
XU$$2035 U$$2035/A U$$2047/B VGND VGND VPWR VPWR U$$2035/X sky130_fd_sc_hd__xor2_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2046 U$$4512/A1 U$$2046/A2 U$$4514/A1 U$$2046/B2 VGND VGND VPWR VPWR U$$2047/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1301 U$$342/A1 U$$1323/A2 U$$70/A1 U$$1307/B2 VGND VGND VPWR VPWR U$$1302/A sky130_fd_sc_hd__a22o_1
XU$$1312 U$$1312/A U$$1316/B VGND VGND VPWR VPWR U$$1312/X sky130_fd_sc_hd__xor2_1
XU$$2057 U$$2178/B VGND VGND VPWR VPWR U$$2057/Y sky130_fd_sc_hd__inv_1
XFILLER_188_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1323 U$$2282/A1 U$$1323/A2 U$$92/A1 U$$1349/B2 VGND VGND VPWR VPWR U$$1324/A sky130_fd_sc_hd__a22o_1
XU$$2068 U$$2068/A U$$2100/B VGND VGND VPWR VPWR U$$2068/X sky130_fd_sc_hd__xor2_1
XU$$1334 U$$1334/A U$$1338/B VGND VGND VPWR VPWR U$$1334/X sky130_fd_sc_hd__xor2_1
XU$$2079 U$$2625/B1 U$$2093/A2 U$$2492/A1 U$$2093/B2 VGND VGND VPWR VPWR U$$2080/A
+ sky130_fd_sc_hd__a22o_1
XU$$1345 U$$932/B1 U$$1367/A2 U$$799/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1346/A sky130_fd_sc_hd__a22o_1
XFILLER_206_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1356 U$$1356/A U$$1366/B VGND VGND VPWR VPWR U$$1356/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_114_1 U$$3826/X U$$3959/X VGND VGND VPWR VPWR dadda_fa_4_115_2/B dadda_ha_3_114_1/SUM
+ sky130_fd_sc_hd__ha_1
XU$$1367 U$$1504/A1 U$$1367/A2 U$$1367/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1368/A
+ sky130_fd_sc_hd__a22o_1
XU$$1378 U$$1515/A1 U$$1448/A2 U$$969/A1 U$$1448/B2 VGND VGND VPWR VPWR U$$1379/A
+ sky130_fd_sc_hd__a22o_1
XU$$1389 U$$1389/A U$$1399/B VGND VGND VPWR VPWR U$$1389/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_106_0 dadda_fa_7_106_0/A dadda_fa_7_106_0/B dadda_fa_7_106_0/CIN VGND
+ VGND VPWR VPWR _403_/D _274_/D sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_10_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _342_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1150 final_adder.U$$899/A1 final_adder.U$$837/X VGND VGND VPWR VPWR
+ output286/A sky130_fd_sc_hd__xor2_2
XFILLER_156_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_988 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_51_0 input203/X dadda_fa_2_51_0/B dadda_fa_2_51_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_52_0/B dadda_fa_3_51_2/B sky130_fd_sc_hd__fa_1
XFILLER_61_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$30 _326_/Q _198_/Q VGND VGND VPWR VPWR final_adder.U$$995/B1 final_adder.U$$224/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$41 _337_/Q _209_/Q VGND VGND VPWR VPWR final_adder.U$$215/B1 final_adder.U$$214/B
+ sky130_fd_sc_hd__ha_1
XFILLER_80_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3270 U$$3270/A U$$3287/A VGND VGND VPWR VPWR U$$3270/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$52 _348_/Q _220_/Q VGND VGND VPWR VPWR final_adder.U$$973/B1 final_adder.U$$202/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3281 U$$3281/A1 U$$3285/A2 U$$3281/B1 U$$3285/B2 VGND VGND VPWR VPWR U$$3282/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$63 _359_/Q _231_/Q VGND VGND VPWR VPWR final_adder.U$$193/B1 final_adder.U$$192/B
+ sky130_fd_sc_hd__ha_1
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3292 U$$3290/Y input43/X U$$3288/A U$$3291/X U$$3288/Y VGND VGND VPWR VPWR U$$3292/X
+ sky130_fd_sc_hd__a32o_4
Xfinal_adder.U$$74 _370_/Q _242_/Q VGND VGND VPWR VPWR final_adder.U$$951/B1 final_adder.U$$180/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$85 _381_/Q _253_/Q VGND VGND VPWR VPWR final_adder.U$$171/B1 final_adder.U$$170/B
+ sky130_fd_sc_hd__ha_1
XFILLER_110_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$96 _392_/Q _264_/Q VGND VGND VPWR VPWR final_adder.U$$929/B1 final_adder.U$$158/A
+ sky130_fd_sc_hd__ha_1
XU$$2580 U$$2717/A1 U$$2588/A2 U$$4500/A1 U$$2588/B2 VGND VGND VPWR VPWR U$$2581/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2591 U$$2591/A U$$2602/A VGND VGND VPWR VPWR U$$2591/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1890 U$$1890/A U$$1917/A VGND VGND VPWR VPWR U$$1890/X sky130_fd_sc_hd__xor2_1
XFILLER_142_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_80_2 dadda_fa_4_80_2/A dadda_fa_4_80_2/B dadda_fa_4_80_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_81_0/CIN dadda_fa_5_80_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_162_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_73_1 dadda_fa_4_73_1/A dadda_fa_4_73_1/B dadda_fa_4_73_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/B dadda_fa_5_73_1/B sky130_fd_sc_hd__fa_1
XFILLER_150_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_89_1 U$$2180/X U$$2313/X U$$2446/X VGND VGND VPWR VPWR dadda_fa_2_90_4/A
+ dadda_fa_2_89_5/B sky130_fd_sc_hd__fa_1
XFILLER_116_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_50_0 dadda_fa_7_50_0/A dadda_fa_7_50_0/B dadda_fa_7_50_0/CIN VGND VGND
+ VPWR VPWR _347_/D _218_/D sky130_fd_sc_hd__fa_2
XFILLER_118_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_66_0 dadda_fa_4_66_0/A dadda_fa_4_66_0/B dadda_fa_4_66_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/A dadda_fa_5_66_1/A sky130_fd_sc_hd__fa_1
XTAP_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$520 final_adder.U$$528/B final_adder.U$$520/B VGND VGND VPWR VPWR
+ final_adder.U$$640/B sky130_fd_sc_hd__and2_1
XTAP_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$531 final_adder.U$$530/B final_adder.U$$415/X final_adder.U$$407/X
+ VGND VGND VPWR VPWR final_adder.U$$531/X sky130_fd_sc_hd__a21o_1
XTAP_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$542 final_adder.U$$550/B final_adder.U$$542/B VGND VGND VPWR VPWR
+ final_adder.U$$662/B sky130_fd_sc_hd__and2_1
XTAP_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$553 final_adder.U$$552/B final_adder.U$$437/X final_adder.U$$429/X
+ VGND VGND VPWR VPWR final_adder.U$$553/X sky130_fd_sc_hd__a21o_1
XTAP_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$564 final_adder.U$$572/B final_adder.U$$564/B VGND VGND VPWR VPWR
+ final_adder.U$$684/B sky130_fd_sc_hd__and2_1
XFILLER_151_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$403 U$$403/A U$$411/A VGND VGND VPWR VPWR U$$403/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$575 final_adder.U$$574/B final_adder.U$$459/X final_adder.U$$451/X
+ VGND VGND VPWR VPWR final_adder.U$$575/X sky130_fd_sc_hd__a21o_1
XTAP_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$414 U$$546/B U$$414/B VGND VGND VPWR VPWR U$$414/X sky130_fd_sc_hd__and2_1
XFILLER_72_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$586 final_adder.U$$594/B final_adder.U$$586/B VGND VGND VPWR VPWR
+ final_adder.U$$706/B sky130_fd_sc_hd__and2_1
XU$$425 U$$836/A1 U$$437/A2 U$$16/A1 U$$437/B2 VGND VGND VPWR VPWR U$$426/A sky130_fd_sc_hd__a22o_1
XTAP_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater790 U$$2608/X VGND VGND VPWR VPWR U$$2711/B2 sky130_fd_sc_hd__buf_6
XFILLER_205_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$597 final_adder.U$$596/B final_adder.U$$481/X final_adder.U$$473/X
+ VGND VGND VPWR VPWR final_adder.U$$597/X sky130_fd_sc_hd__a21o_1
XU$$436 U$$436/A U$$436/B VGND VGND VPWR VPWR U$$436/X sky130_fd_sc_hd__xor2_1
XTAP_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$447 U$$36/A1 U$$473/A2 U$$38/A1 U$$473/B2 VGND VGND VPWR VPWR U$$448/A sky130_fd_sc_hd__a22o_1
XFILLER_189_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$458 U$$458/A U$$492/B VGND VGND VPWR VPWR U$$458/X sky130_fd_sc_hd__xor2_1
XU$$469 U$$878/B1 U$$473/A2 U$$745/A1 U$$473/B2 VGND VGND VPWR VPWR U$$470/A sky130_fd_sc_hd__a22o_1
XFILLER_189_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1303 U$$3349/B VGND VGND VPWR VPWR U$$3321/B sky130_fd_sc_hd__buf_8
XFILLER_126_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1314 U$$3244/B VGND VGND VPWR VPWR U$$3242/B sky130_fd_sc_hd__buf_8
XFILLER_176_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1325 U$$3133/B VGND VGND VPWR VPWR U$$3125/B sky130_fd_sc_hd__buf_12
XFILLER_154_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1336 U$$3008/B VGND VGND VPWR VPWR U$$2996/B sky130_fd_sc_hd__buf_6
XFILLER_5_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1347 U$$2845/B VGND VGND VPWR VPWR U$$2837/B sky130_fd_sc_hd__buf_6
XFILLER_126_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1358 U$$2658/B VGND VGND VPWR VPWR U$$2650/B sky130_fd_sc_hd__buf_6
XFILLER_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1369 U$$2525/B VGND VGND VPWR VPWR U$$2491/B sky130_fd_sc_hd__buf_6
XFILLER_84_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_830 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_59_clk _219_/CLK VGND VGND VPWR VPWR _211_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_471 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$970 U$$970/A U$$980/B VGND VGND VPWR VPWR U$$970/X sky130_fd_sc_hd__xor2_1
XFILLER_35_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1120 U$$1666/B1 U$$1136/A2 U$$985/A1 U$$1136/B2 VGND VGND VPWR VPWR U$$1121/A
+ sky130_fd_sc_hd__a22o_1
XU$$981 U$$981/A1 U$$999/A2 U$$983/A1 U$$999/B2 VGND VGND VPWR VPWR U$$982/A sky130_fd_sc_hd__a22o_1
XFILLER_211_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$992 U$$992/A U$$994/B VGND VGND VPWR VPWR U$$992/X sky130_fd_sc_hd__xor2_1
XU$$1131 U$$1131/A U$$1187/B VGND VGND VPWR VPWR U$$1131/X sky130_fd_sc_hd__xor2_1
XU$$1142 U$$731/A1 U$$1190/A2 U$$733/A1 U$$1190/B2 VGND VGND VPWR VPWR U$$1143/A sky130_fd_sc_hd__a22o_1
XU$$1153 U$$1153/A U$$1195/B VGND VGND VPWR VPWR U$$1153/X sky130_fd_sc_hd__xor2_1
XFILLER_50_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1164 U$$2123/A1 U$$1190/A2 U$$616/B1 U$$1190/B2 VGND VGND VPWR VPWR U$$1165/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1175 U$$1175/A U$$1175/B VGND VGND VPWR VPWR U$$1175/X sky130_fd_sc_hd__xor2_1
XFILLER_31_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1186 U$$773/B1 U$$1190/A2 U$$640/A1 U$$1190/B2 VGND VGND VPWR VPWR U$$1187/A sky130_fd_sc_hd__a22o_1
XFILLER_148_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1197 U$$1197/A U$$1205/B VGND VGND VPWR VPWR U$$1197/X sky130_fd_sc_hd__xor2_1
XFILLER_203_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_90_1 dadda_fa_5_90_1/A dadda_fa_5_90_1/B dadda_fa_5_90_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_91_0/B dadda_fa_7_90_0/A sky130_fd_sc_hd__fa_1
XFILLER_191_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_83_0 dadda_fa_5_83_0/A dadda_fa_5_83_0/B dadda_fa_5_83_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_84_0/A dadda_fa_6_83_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_172_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_99_0 U$$2465/Y U$$2599/X U$$2732/X VGND VGND VPWR VPWR dadda_fa_3_100_1/A
+ dadda_fa_3_99_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_75_7 U$$4413/X input229/X dadda_fa_1_75_7/CIN VGND VGND VPWR VPWR dadda_fa_2_76_2/CIN
+ dadda_fa_2_75_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_112_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_68_6 dadda_fa_1_68_6/A dadda_fa_1_68_6/B dadda_fa_1_68_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_2/B dadda_fa_2_68_5/B sky130_fd_sc_hd__fa_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_814 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 _386_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$545_1837 VGND VGND VPWR VPWR U$$545_1837/HI U$$545/B1 sky130_fd_sc_hd__conb_1
XFILLER_96_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_474 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_98_0 dadda_fa_7_98_0/A dadda_fa_7_98_0/B dadda_fa_7_98_0/CIN VGND VGND
+ VPWR VPWR _395_/D _266_/D sky130_fd_sc_hd__fa_1
XFILLER_167_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3431_1749 VGND VGND VPWR VPWR U$$3431_1749/HI U$$3431/A1 sky130_fd_sc_hd__conb_1
XFILLER_136_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_113_0 dadda_fa_6_113_0/A dadda_fa_6_113_0/B dadda_fa_6_113_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_114_0/B dadda_fa_7_113_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$350 final_adder.U$$352/B final_adder.U$$350/B VGND VGND VPWR VPWR
+ final_adder.U$$476/B sky130_fd_sc_hd__and2_1
XTAP_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$361 final_adder.U$$360/B final_adder.U$$235/X final_adder.U$$233/X
+ VGND VGND VPWR VPWR final_adder.U$$361/X sky130_fd_sc_hd__a21o_1
XTAP_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$200 U$$200/A U$$218/B VGND VGND VPWR VPWR U$$200/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$372 final_adder.U$$374/B final_adder.U$$372/B VGND VGND VPWR VPWR
+ final_adder.U$$498/B sky130_fd_sc_hd__and2_1
XTAP_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$211 U$$74/A1 U$$259/A2 U$$76/A1 U$$259/B2 VGND VGND VPWR VPWR U$$212/A sky130_fd_sc_hd__a22o_1
XTAP_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$222 U$$222/A U$$264/B VGND VGND VPWR VPWR U$$222/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_33_3 dadda_fa_3_33_3/A dadda_fa_3_33_3/B dadda_fa_3_33_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_34_1/B dadda_fa_4_33_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$394 final_adder.U$$398/B final_adder.U$$394/B VGND VGND VPWR VPWR
+ final_adder.U$$518/B sky130_fd_sc_hd__and2_1
XTAP_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$233 U$$916/B1 U$$259/A2 U$$98/A1 U$$259/B2 VGND VGND VPWR VPWR U$$234/A sky130_fd_sc_hd__a22o_1
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$244 U$$244/A U$$244/B VGND VGND VPWR VPWR U$$244/X sky130_fd_sc_hd__xor2_1
XTAP_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$255 U$$392/A1 U$$257/A2 U$$942/A1 U$$257/B2 VGND VGND VPWR VPWR U$$256/A sky130_fd_sc_hd__a22o_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$266 U$$266/A U$$272/B VGND VGND VPWR VPWR U$$266/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_26_2 U$$1820/B input175/X dadda_fa_3_26_2/CIN VGND VGND VPWR VPWR dadda_fa_4_27_1/A
+ dadda_fa_4_26_2/B sky130_fd_sc_hd__fa_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$277 U$$411/A U$$277/B VGND VGND VPWR VPWR U$$277/X sky130_fd_sc_hd__and2_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$288 U$$14/A1 U$$316/A2 U$$16/A1 U$$316/B2 VGND VGND VPWR VPWR U$$289/A sky130_fd_sc_hd__a22o_1
XFILLER_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$299 U$$299/A U$$379/B VGND VGND VPWR VPWR U$$299/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_3_19_1 U$$444/X U$$577/X U$$710/X VGND VGND VPWR VPWR dadda_fa_4_20_1/A
+ dadda_fa_4_19_2/B sky130_fd_sc_hd__fa_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$5 U$$3/B U$$5/A2 U$$1/A U$$0/Y VGND VGND VPWR VPWR U$$5/X sky130_fd_sc_hd__a22o_1
XFILLER_126_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1100 U$$2202/A1 VGND VGND VPWR VPWR U$$2063/B1 sky130_fd_sc_hd__buf_6
XFILLER_154_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1111 U$$3880/B1 VGND VGND VPWR VPWR U$$44/B1 sky130_fd_sc_hd__buf_6
XFILLER_126_443 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput308 output308/A VGND VGND VPWR VPWR o[30] sky130_fd_sc_hd__buf_2
XFILLER_142_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1122 U$$179/A1 VGND VGND VPWR VPWR U$$42/A1 sky130_fd_sc_hd__buf_4
Xoutput319 output319/A VGND VGND VPWR VPWR o[40] sky130_fd_sc_hd__buf_2
XFILLER_142_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1133 U$$4011/B1 VGND VGND VPWR VPWR U$$997/B1 sky130_fd_sc_hd__buf_6
Xrepeater1144 U$$4422/A1 VGND VGND VPWR VPWR U$$3737/A1 sky130_fd_sc_hd__buf_8
Xrepeater1155 U$$998/B VGND VGND VPWR VPWR U$$996/B sky130_fd_sc_hd__buf_6
XFILLER_142_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1166 U$$3183/B1 VGND VGND VPWR VPWR U$$2363/A1 sky130_fd_sc_hd__buf_6
Xrepeater1177 U$$32/A1 VGND VGND VPWR VPWR U$$717/A1 sky130_fd_sc_hd__clkbuf_4
Xrepeater1188 input66/X VGND VGND VPWR VPWR U$$28/A1 sky130_fd_sc_hd__buf_4
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1199 U$$1515/A1 VGND VGND VPWR VPWR U$$2198/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_2_78_5 dadda_fa_2_78_5/A dadda_fa_2_78_5/B dadda_fa_2_78_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_79_2/A dadda_fa_4_78_0/A sky130_fd_sc_hd__fa_2
XFILLER_68_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_108_1 dadda_fa_5_108_1/A dadda_fa_5_108_1/B dadda_fa_5_108_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_109_0/B dadda_fa_7_108_0/A sky130_fd_sc_hd__fa_1
XFILLER_118_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_80_5 U$$3093/X U$$3226/X U$$3359/X VGND VGND VPWR VPWR dadda_fa_2_81_2/B
+ dadda_fa_2_80_5/A sky130_fd_sc_hd__fa_1
XFILLER_120_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_73_4 U$$3478/X U$$3611/X U$$3744/X VGND VGND VPWR VPWR dadda_fa_2_74_1/CIN
+ dadda_fa_2_73_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_66_3 U$$3730/X U$$3863/X U$$3996/X VGND VGND VPWR VPWR dadda_fa_2_67_1/B
+ dadda_fa_2_66_4/B sky130_fd_sc_hd__fa_1
XFILLER_100_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_43_2 dadda_fa_4_43_2/A dadda_fa_4_43_2/B dadda_fa_4_43_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_44_0/CIN dadda_fa_5_43_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_59_2 U$$2386/X U$$2519/X U$$2652/X VGND VGND VPWR VPWR dadda_fa_2_60_1/A
+ dadda_fa_2_59_4/A sky130_fd_sc_hd__fa_1
XFILLER_100_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_36_1 dadda_fa_4_36_1/A dadda_fa_4_36_1/B dadda_fa_4_36_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/B dadda_fa_5_36_1/B sky130_fd_sc_hd__fa_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_13_0 dadda_fa_7_13_0/A dadda_fa_7_13_0/B dadda_fa_7_13_0/CIN VGND VGND
+ VPWR VPWR _310_/D _181_/D sky130_fd_sc_hd__fa_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_29_0 dadda_fa_4_29_0/A dadda_fa_4_29_0/B dadda_fa_4_29_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/A dadda_fa_5_29_1/A sky130_fd_sc_hd__fa_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_260_ _414_/CLK _260_/D VGND VGND VPWR VPWR _260_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_191_ _326_/CLK _191_/D VGND VGND VPWR VPWR _191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1056 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4504 U$$4504/A1 U$$4388/X U$$4506/A1 U$$4512/B2 VGND VGND VPWR VPWR U$$4505/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4515 U$$4515/A U$$4515/B VGND VGND VPWR VPWR U$$4515/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_0_61_2 U$$927/X U$$1060/X U$$1193/X VGND VGND VPWR VPWR dadda_fa_1_62_6/B
+ dadda_fa_1_61_8/B sky130_fd_sc_hd__fa_1
XFILLER_49_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3803 input107/X U$$3819/A2 input108/X U$$3819/B2 VGND VGND VPWR VPWR U$$3804/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3814 U$$3814/A U$$3814/B VGND VGND VPWR VPWR U$$3814/X sky130_fd_sc_hd__xor2_1
XU$$18 U$$18/A1 U$$42/A2 U$$20/A1 U$$42/B2 VGND VGND VPWR VPWR U$$19/A sky130_fd_sc_hd__a22o_1
XTAP_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$29 U$$29/A U$$51/B VGND VGND VPWR VPWR U$$29/X sky130_fd_sc_hd__xor2_1
XTAP_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3825 U$$3960/B1 U$$3833/A2 U$$4099/B1 U$$3833/B2 VGND VGND VPWR VPWR U$$3826/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3836 U$$3836/A VGND VGND VPWR VPWR U$$3836/Y sky130_fd_sc_hd__inv_1
XTAP_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_31_0 U$$1931/X U$$2064/X input181/X VGND VGND VPWR VPWR dadda_fa_4_32_0/B
+ dadda_fa_4_31_1/CIN sky130_fd_sc_hd__fa_1
XU$$3847 U$$3847/A U$$3879/B VGND VGND VPWR VPWR U$$3847/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$180 final_adder.U$$180/A final_adder.U$$180/B VGND VGND VPWR VPWR
+ final_adder.U$$308/B sky130_fd_sc_hd__and2_1
XFILLER_166_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3858 U$$4269/A1 U$$3874/A2 U$$4269/B1 U$$3874/B2 VGND VGND VPWR VPWR U$$3859/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$191 final_adder.U$$190/B final_adder.U$$961/B1 final_adder.U$$191/B1
+ VGND VGND VPWR VPWR final_adder.U$$191/X sky130_fd_sc_hd__a21o_1
XTAP_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3869 U$$3869/A U$$3903/B VGND VGND VPWR VPWR U$$3869/X sky130_fd_sc_hd__xor2_1
XFILLER_79_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_389_ _414_/CLK _389_/D VGND VGND VPWR VPWR _389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_90_4 dadda_fa_2_90_4/A dadda_fa_2_90_4/B dadda_fa_2_90_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_91_1/CIN dadda_fa_3_90_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_56_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_83_3 dadda_fa_2_83_3/A dadda_fa_2_83_3/B dadda_fa_2_83_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/B dadda_fa_3_83_3/B sky130_fd_sc_hd__fa_1
XFILLER_181_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_76_2 dadda_fa_2_76_2/A dadda_fa_2_76_2/B dadda_fa_2_76_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/A dadda_fa_3_76_3/A sky130_fd_sc_hd__fa_1
Xdadda_fa_5_53_1 dadda_fa_5_53_1/A dadda_fa_5_53_1/B dadda_fa_5_53_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_54_0/B dadda_fa_7_53_0/A sky130_fd_sc_hd__fa_1
Xdadda_fa_2_69_1 dadda_fa_2_69_1/A dadda_fa_2_69_1/B dadda_fa_2_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_0/CIN dadda_fa_3_69_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_842 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_46_0 dadda_fa_5_46_0/A dadda_fa_5_46_0/B dadda_fa_5_46_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_47_0/A dadda_fa_6_46_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_120_0 U$$4503/X input152/X dadda_fa_5_120_0/CIN VGND VGND VPWR VPWR dadda_fa_6_121_0/A
+ dadda_fa_6_120_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_30_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_71_1 U$$2543/X U$$2676/X U$$2809/X VGND VGND VPWR VPWR dadda_fa_2_72_0/CIN
+ dadda_fa_2_71_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_120_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_64_0 U$$2529/X U$$2662/X U$$2795/X VGND VGND VPWR VPWR dadda_fa_2_65_0/B
+ dadda_fa_2_64_3/B sky130_fd_sc_hd__fa_1
XFILLER_8_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_396 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2409 U$$2957/A1 U$$2435/A2 U$$2409/B1 U$$2435/B2 VGND VGND VPWR VPWR U$$2410/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1708 U$$3215/A1 U$$1750/A2 U$$1984/A1 U$$1750/B2 VGND VGND VPWR VPWR U$$1709/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1719 U$$1719/A U$$1721/B VGND VGND VPWR VPWR U$$1719/X sky130_fd_sc_hd__xor2_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_312_ _314_/CLK _312_/D VGND VGND VPWR VPWR _312_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_499 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_243_ _373_/CLK _243_/D VGND VGND VPWR VPWR _243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_1014 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput18 a[25] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__buf_6
X_174_ _304_/CLK _174_/D VGND VGND VPWR VPWR _174_/Q sky130_fd_sc_hd__dfxtp_1
Xinput29 a[35] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_868 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_93_2 dadda_fa_3_93_2/A dadda_fa_3_93_2/B dadda_fa_3_93_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_1/A dadda_fa_4_93_2/B sky130_fd_sc_hd__fa_1
XFILLER_202_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_86_1 dadda_fa_3_86_1/A dadda_fa_3_86_1/B dadda_fa_3_86_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_0/CIN dadda_fa_4_86_2/A sky130_fd_sc_hd__fa_1
XFILLER_184_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_63_0 dadda_fa_6_63_0/A dadda_fa_6_63_0/B dadda_fa_6_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_64_0/B dadda_fa_7_63_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_79_0 dadda_fa_3_79_0/A dadda_fa_3_79_0/B dadda_fa_3_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_0/B dadda_fa_4_79_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_ha_0_53_0 U$$113/X U$$246/X VGND VGND VPWR VPWR dadda_fa_1_54_8/B dadda_fa_2_53_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_111_416 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater608 U$$263/A2 VGND VGND VPWR VPWR U$$217/A2 sky130_fd_sc_hd__buf_6
XU$$4301 U$$4438/A1 U$$4381/A2 U$$4440/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4302/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater619 U$$1470/A2 VGND VGND VPWR VPWR U$$1422/A2 sky130_fd_sc_hd__buf_4
XU$$4312 U$$4312/A U$$4370/B VGND VGND VPWR VPWR U$$4312/X sky130_fd_sc_hd__xor2_1
XFILLER_42_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4323 U$$4460/A1 U$$4327/A2 U$$4323/B1 U$$4327/B2 VGND VGND VPWR VPWR U$$4324/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4334 U$$4334/A U$$4354/B VGND VGND VPWR VPWR U$$4334/X sky130_fd_sc_hd__xor2_1
XU$$4345 U$$783/A1 U$$4361/A2 U$$4484/A1 U$$4361/B2 VGND VGND VPWR VPWR U$$4346/A
+ sky130_fd_sc_hd__a22o_1
XU$$3600 U$$3737/A1 U$$3636/A2 U$$3737/B1 U$$3636/B2 VGND VGND VPWR VPWR U$$3601/A
+ sky130_fd_sc_hd__a22o_1
XU$$4356 U$$4356/A U$$4366/B VGND VGND VPWR VPWR U$$4356/X sky130_fd_sc_hd__xor2_1
XFILLER_133_1198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3611 U$$3611/A U$$3697/B VGND VGND VPWR VPWR U$$3611/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_115_1 U$$4360/X U$$4493/X input146/X VGND VGND VPWR VPWR dadda_fa_5_116_0/B
+ dadda_fa_5_115_1/B sky130_fd_sc_hd__fa_1
XU$$3622 input83/X U$$3644/A2 U$$3761/A1 U$$3644/B2 VGND VGND VPWR VPWR U$$3623/A
+ sky130_fd_sc_hd__a22o_1
XU$$4367 U$$4504/A1 U$$4369/A2 U$$4506/A1 U$$4369/B2 VGND VGND VPWR VPWR U$$4368/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3633 U$$3633/A U$$3637/B VGND VGND VPWR VPWR U$$3633/X sky130_fd_sc_hd__xor2_1
XFILLER_53_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4378 U$$4378/A U$$4382/B VGND VGND VPWR VPWR U$$4378/X sky130_fd_sc_hd__xor2_1
XFILLER_92_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4389 U$$4387/B U$$4384/A U$$4389/B1 U$$4384/Y VGND VGND VPWR VPWR U$$4389/X sky130_fd_sc_hd__a22o_4
XFILLER_19_975 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3644 U$$3644/A1 U$$3644/A2 U$$3644/B1 U$$3644/B2 VGND VGND VPWR VPWR U$$3645/A
+ sky130_fd_sc_hd__a22o_1
XU$$2910 U$$2910/A U$$2996/B VGND VGND VPWR VPWR U$$2910/X sky130_fd_sc_hd__xor2_1
XU$$3655 U$$3655/A U$$3665/B VGND VGND VPWR VPWR U$$3655/X sky130_fd_sc_hd__xor2_1
XFILLER_52_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3666 U$$3801/B1 U$$3680/A2 U$$4077/B1 U$$3680/B2 VGND VGND VPWR VPWR U$$3667/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_108_0 dadda_fa_4_108_0/A dadda_fa_4_108_0/B dadda_fa_4_108_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/A dadda_fa_5_108_1/A sky130_fd_sc_hd__fa_1
XU$$2921 U$$3058/A1 U$$2921/A2 U$$3606/B1 U$$2921/B2 VGND VGND VPWR VPWR U$$2922/A
+ sky130_fd_sc_hd__a22o_1
XU$$3677 U$$3677/A U$$3683/B VGND VGND VPWR VPWR U$$3677/X sky130_fd_sc_hd__xor2_1
XU$$2932 U$$2932/A U$$2978/B VGND VGND VPWR VPWR U$$2932/X sky130_fd_sc_hd__xor2_1
XFILLER_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3688 input119/X U$$3696/A2 U$$4099/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3689/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2943 U$$3078/B1 U$$2967/A2 U$$3356/A1 U$$2967/B2 VGND VGND VPWR VPWR U$$2944/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2954 U$$2954/A U$$2996/B VGND VGND VPWR VPWR U$$2954/X sky130_fd_sc_hd__xor2_1
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3699 input49/X VGND VGND VPWR VPWR U$$3699/Y sky130_fd_sc_hd__inv_1
XU$$2965 U$$3376/A1 U$$2977/A2 U$$3378/A1 U$$2979/B2 VGND VGND VPWR VPWR U$$2966/A
+ sky130_fd_sc_hd__a22o_1
XU$$2976 U$$2976/A U$$2978/B VGND VGND VPWR VPWR U$$2976/X sky130_fd_sc_hd__xor2_1
XFILLER_33_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2987 U$$384/A1 U$$2995/A2 U$$521/B1 U$$2995/B2 VGND VGND VPWR VPWR U$$2988/A sky130_fd_sc_hd__a22o_1
XANTENNA_270 U$$1877/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2998 U$$2998/A U$$3013/A VGND VGND VPWR VPWR U$$2998/X sky130_fd_sc_hd__xor2_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_81_0 U$$4425/X input236/X dadda_fa_2_81_0/CIN VGND VGND VPWR VPWR dadda_fa_3_82_0/B
+ dadda_fa_3_81_2/B sky130_fd_sc_hd__fa_1
XFILLER_88_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_1_51_8 U$$3301/X U$$3434/X VGND VGND VPWR VPWR dadda_fa_2_52_3/A dadda_fa_3_51_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_115_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$905 final_adder.U$$134/A final_adder.U$$843/X final_adder.U$$905/B1
+ VGND VGND VPWR VPWR final_adder.U$$905/X sky130_fd_sc_hd__a21o_1
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$927 final_adder.U$$156/A final_adder.U$$865/X final_adder.U$$927/B1
+ VGND VGND VPWR VPWR final_adder.U$$927/X sky130_fd_sc_hd__a21o_1
XFILLER_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$949 final_adder.U$$178/A final_adder.U$$887/X final_adder.U$$949/B1
+ VGND VGND VPWR VPWR final_adder.U$$949/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_1_50_6 U$$2501/X U$$2634/X U$$2767/X VGND VGND VPWR VPWR dadda_fa_2_51_2/B
+ dadda_fa_2_50_5/B sky130_fd_sc_hd__fa_1
XFILLER_68_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_2_0 U$$160/B input179/X dadda_ha_6_2_0/SUM VGND VGND VPWR VPWR _299_/D
+ _170_/D sky130_fd_sc_hd__fa_1
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_775 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_747 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_80_0 dadda_fa_7_80_0/A dadda_fa_7_80_0/B dadda_fa_7_80_0/CIN VGND VGND
+ VPWR VPWR _377_/D _248_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_96_0 dadda_fa_4_96_0/A dadda_fa_4_96_0/B dadda_fa_4_96_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/A dadda_fa_5_96_1/A sky130_fd_sc_hd__fa_1
XFILLER_153_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2206 U$$3300/B1 U$$2226/A2 U$$2206/B1 U$$2226/B2 VGND VGND VPWR VPWR U$$2207/A
+ sky130_fd_sc_hd__a22o_1
XU$$2217 U$$2217/A U$$2273/B VGND VGND VPWR VPWR U$$2217/X sky130_fd_sc_hd__xor2_1
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2228 U$$995/A1 U$$2252/A2 U$$4011/A1 U$$2252/B2 VGND VGND VPWR VPWR U$$2229/A
+ sky130_fd_sc_hd__a22o_1
XU$$4385_1766 VGND VGND VPWR VPWR U$$4385_1766/HI U$$4385/A sky130_fd_sc_hd__conb_1
XU$$2239 U$$2239/A U$$2285/B VGND VGND VPWR VPWR U$$2239/X sky130_fd_sc_hd__xor2_1
XFILLER_43_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1505 U$$1505/A U$$1507/A VGND VGND VPWR VPWR U$$1505/X sky130_fd_sc_hd__xor2_1
XFILLER_103_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1516 U$$1516/A U$$1574/B VGND VGND VPWR VPWR U$$1516/X sky130_fd_sc_hd__xor2_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1527 U$$1799/B1 U$$1545/A2 U$$1666/A1 U$$1545/B2 VGND VGND VPWR VPWR U$$1528/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1538 U$$1538/A U$$1574/B VGND VGND VPWR VPWR U$$1538/X sky130_fd_sc_hd__xor2_1
XFILLER_15_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1549 U$$864/A1 U$$1557/A2 U$$864/B1 U$$1557/B2 VGND VGND VPWR VPWR U$$1550/A sky130_fd_sc_hd__a22o_1
XFILLER_179_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_972 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_226_ _359_/CLK _226_/D VGND VGND VPWR VPWR _226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_839 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_60_5 dadda_fa_2_60_5/A dadda_fa_2_60_5/B dadda_fa_2_60_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_61_2/A dadda_fa_4_60_0/A sky130_fd_sc_hd__fa_2
Xrepeater405 U$$805/A2 VGND VGND VPWR VPWR U$$759/A2 sky130_fd_sc_hd__buf_4
Xrepeater416 U$$4251/X VGND VGND VPWR VPWR U$$4297/A2 sky130_fd_sc_hd__buf_4
Xrepeater427 U$$415/X VGND VGND VPWR VPWR U$$527/A2 sky130_fd_sc_hd__buf_6
XFILLER_65_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_53_4 dadda_fa_2_53_4/A dadda_fa_2_53_4/B dadda_fa_2_53_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_1/CIN dadda_fa_3_53_3/CIN sky130_fd_sc_hd__fa_1
XU$$4120 U$$4394/A1 U$$4144/A2 U$$4396/A1 U$$4144/B2 VGND VGND VPWR VPWR U$$4121/A
+ sky130_fd_sc_hd__a22o_1
Xrepeater438 U$$4114/X VGND VGND VPWR VPWR U$$4240/A2 sky130_fd_sc_hd__buf_4
Xrepeater449 U$$4079/A2 VGND VGND VPWR VPWR U$$4077/A2 sky130_fd_sc_hd__clkbuf_4
XU$$4131 U$$4131/A U$$4246/A VGND VGND VPWR VPWR U$$4131/X sky130_fd_sc_hd__xor2_1
XFILLER_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4142 U$$4277/B1 U$$4144/A2 U$$4144/A1 U$$4144/B2 VGND VGND VPWR VPWR U$$4143/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_46_3 dadda_fa_2_46_3/A dadda_fa_2_46_3/B dadda_fa_2_46_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/B dadda_fa_3_46_3/B sky130_fd_sc_hd__fa_1
XU$$4153 U$$4153/A U$$4189/B VGND VGND VPWR VPWR U$$4153/X sky130_fd_sc_hd__xor2_1
XFILLER_38_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4164 U$$4438/A1 U$$4164/A2 U$$4440/A1 U$$4164/B2 VGND VGND VPWR VPWR U$$4165/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4175 U$$4175/A U$$4246/A VGND VGND VPWR VPWR U$$4175/X sky130_fd_sc_hd__xor2_1
XU$$3430 U$$3428/B U$$3377/B input46/X U$$3425/Y VGND VGND VPWR VPWR U$$3430/X sky130_fd_sc_hd__a22o_4
XU$$3441 U$$3578/A1 U$$3527/A2 U$$3578/B1 U$$3527/B2 VGND VGND VPWR VPWR U$$3442/A
+ sky130_fd_sc_hd__a22o_1
XU$$4186 U$$4460/A1 U$$4188/A2 input93/X U$$4188/B2 VGND VGND VPWR VPWR U$$4187/A
+ sky130_fd_sc_hd__a22o_1
XU$$4197 U$$4197/A U$$4211/B VGND VGND VPWR VPWR U$$4197/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3452 U$$3452/A U$$3454/B VGND VGND VPWR VPWR U$$3452/X sky130_fd_sc_hd__xor2_1
XU$$3463 U$$3737/A1 U$$3503/A2 U$$3737/B1 U$$3503/B2 VGND VGND VPWR VPWR U$$3464/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_39_2 U$$1947/X U$$2080/X U$$2213/X VGND VGND VPWR VPWR dadda_fa_3_40_1/A
+ dadda_fa_3_39_3/A sky130_fd_sc_hd__fa_1
XFILLER_129_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3474 U$$3474/A U$$3480/B VGND VGND VPWR VPWR U$$3474/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_16_1 dadda_fa_5_16_1/A dadda_fa_5_16_1/B dadda_fa_5_16_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_17_0/B dadda_fa_7_16_0/A sky130_fd_sc_hd__fa_1
XU$$3485 U$$3485/A1 U$$3489/A2 input84/X U$$3489/B2 VGND VGND VPWR VPWR U$$3486/A
+ sky130_fd_sc_hd__a22o_1
XU$$2740 input33/X VGND VGND VPWR VPWR U$$2740/Y sky130_fd_sc_hd__inv_1
XFILLER_94_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2751 U$$2751/A U$$2755/B VGND VGND VPWR VPWR U$$2751/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3496 U$$3496/A U$$3510/B VGND VGND VPWR VPWR U$$3496/X sky130_fd_sc_hd__xor2_1
XFILLER_179_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2762 U$$3447/A1 U$$2782/A2 U$$3584/B1 U$$2782/B2 VGND VGND VPWR VPWR U$$2763/A
+ sky130_fd_sc_hd__a22o_1
XU$$2773 U$$2773/A U$$2783/B VGND VGND VPWR VPWR U$$2773/X sky130_fd_sc_hd__xor2_1
XFILLER_22_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2784 U$$3058/A1 U$$2828/A2 U$$3880/B1 U$$2828/B2 VGND VGND VPWR VPWR U$$2785/A
+ sky130_fd_sc_hd__a22o_1
XU$$2795 U$$2795/A U$$2797/B VGND VGND VPWR VPWR U$$2795/X sky130_fd_sc_hd__xor2_1
XFILLER_21_425 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_1_42_4 U$$1687/X U$$1820/X VGND VGND VPWR VPWR dadda_fa_2_43_4/B dadda_fa_3_42_0/A
+ sky130_fd_sc_hd__ha_1
Xinput208 c[56] VGND VGND VPWR VPWR input208/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput219 c[66] VGND VGND VPWR VPWR input219/X sky130_fd_sc_hd__clkbuf_1
XTAP_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$702 final_adder.U$$718/B final_adder.U$$702/B VGND VGND VPWR VPWR
+ final_adder.U$$782/A sky130_fd_sc_hd__and2_1
XTAP_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$713 final_adder.U$$712/B final_adder.U$$609/X final_adder.U$$593/X
+ VGND VGND VPWR VPWR final_adder.U$$713/X sky130_fd_sc_hd__a21o_1
XTAP_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_4_12_2 U$$829/X U$$919/B VGND VGND VPWR VPWR dadda_fa_5_13_0/CIN dadda_ha_4_12_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_68_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$735 final_adder.U$$718/A final_adder.U$$381/X final_adder.U$$615/X
+ VGND VGND VPWR VPWR final_adder.U$$735/X sky130_fd_sc_hd__a21o_2
XFILLER_84_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$746 final_adder.U$$778/B final_adder.U$$746/B VGND VGND VPWR VPWR
+ final_adder.U$$746/X sky130_fd_sc_hd__and2_1
Xrepeater950 input94/X VGND VGND VPWR VPWR U$$4464/A1 sky130_fd_sc_hd__buf_6
XFILLER_56_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$757 final_adder.U$$756/B final_adder.U$$677/X final_adder.U$$645/X
+ VGND VGND VPWR VPWR final_adder.U$$757/X sky130_fd_sc_hd__a21o_1
Xrepeater961 U$$4460/A1 VGND VGND VPWR VPWR U$$2951/B1 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$768 final_adder.U$$800/B final_adder.U$$768/B VGND VGND VPWR VPWR
+ final_adder.U$$768/X sky130_fd_sc_hd__and2_1
Xrepeater972 U$$4458/A1 VGND VGND VPWR VPWR U$$3088/A1 sky130_fd_sc_hd__buf_6
XFILLER_17_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$607 U$$607/A U$$607/B VGND VGND VPWR VPWR U$$607/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$779 final_adder.U$$778/B final_adder.U$$699/X final_adder.U$$667/X
+ VGND VGND VPWR VPWR final_adder.U$$779/X sky130_fd_sc_hd__a21o_1
XU$$618 U$$892/A1 U$$624/A2 U$$757/A1 U$$624/B2 VGND VGND VPWR VPWR U$$619/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_1_41_2 U$$887/X U$$1020/X U$$1153/X VGND VGND VPWR VPWR dadda_fa_2_42_4/A
+ dadda_fa_2_41_5/CIN sky130_fd_sc_hd__fa_1
Xrepeater983 U$$1187/B VGND VGND VPWR VPWR U$$1137/B sky130_fd_sc_hd__clkbuf_8
XFILLER_99_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater994 U$$4454/A1 VGND VGND VPWR VPWR U$$1714/A1 sky130_fd_sc_hd__buf_4
XU$$629 U$$629/A U$$673/B VGND VGND VPWR VPWR U$$629/X sky130_fd_sc_hd__xor2_1
XFILLER_56_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_1199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_11_0 U$$29/X U$$162/X U$$295/X VGND VGND VPWR VPWR dadda_fa_5_12_0/B dadda_fa_5_11_1/B
+ sky130_fd_sc_hd__fa_1
XFILLER_13_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_90_0_1857 VGND VGND VPWR VPWR dadda_fa_1_90_0/A dadda_fa_1_90_0_1857/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1507 U$$952/A1 VGND VGND VPWR VPWR U$$950/B1 sky130_fd_sc_hd__buf_4
Xrepeater1518 input121/X VGND VGND VPWR VPWR U$$3416/A1 sky130_fd_sc_hd__buf_4
XFILLER_165_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_115_0 U$$3561/Y U$$3695/X U$$3828/X VGND VGND VPWR VPWR dadda_fa_4_116_2/B
+ dadda_fa_4_115_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater1529 U$$99/B VGND VGND VPWR VPWR U$$85/B sky130_fd_sc_hd__buf_8
XFILLER_153_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_63_3 dadda_fa_3_63_3/A dadda_fa_3_63_3/B dadda_fa_3_63_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_64_1/B dadda_fa_4_63_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_58_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_56_2 dadda_fa_3_56_2/A dadda_fa_3_56_2/B dadda_fa_3_56_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_1/A dadda_fa_4_56_2/B sky130_fd_sc_hd__fa_1
XFILLER_58_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_49_1 dadda_fa_3_49_1/A dadda_fa_3_49_1/B dadda_fa_3_49_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_0/CIN dadda_fa_4_49_2/A sky130_fd_sc_hd__fa_1
XFILLER_43_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_26_0 dadda_fa_6_26_0/A dadda_fa_6_26_0/B dadda_fa_6_26_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_27_0/B dadda_fa_7_26_0/CIN sky130_fd_sc_hd__fa_1
XU$$2003 U$$2003/A U$$2043/B VGND VGND VPWR VPWR U$$2003/X sky130_fd_sc_hd__xor2_1
XFILLER_35_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2014 U$$2425/A1 U$$2022/A2 U$$2016/A1 U$$2022/B2 VGND VGND VPWR VPWR U$$2015/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2025 U$$2025/A U$$2054/A VGND VGND VPWR VPWR U$$2025/X sky130_fd_sc_hd__xor2_1
XU$$2036 U$$2445/B1 U$$2046/A2 U$$2312/A1 U$$2046/B2 VGND VGND VPWR VPWR U$$2037/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2047 U$$2047/A U$$2047/B VGND VGND VPWR VPWR U$$2047/X sky130_fd_sc_hd__xor2_1
XU$$1302 U$$1302/A U$$1354/B VGND VGND VPWR VPWR U$$1302/X sky130_fd_sc_hd__xor2_1
XU$$1313 U$$902/A1 U$$1361/A2 U$$4055/A1 U$$1355/B2 VGND VGND VPWR VPWR U$$1314/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2058 input25/X U$$2058/B VGND VGND VPWR VPWR U$$2058/X sky130_fd_sc_hd__and2_1
XU$$1324 U$$1324/A U$$1354/B VGND VGND VPWR VPWR U$$1324/X sky130_fd_sc_hd__xor2_1
XU$$2069 U$$2069/A1 U$$2099/A2 U$$2206/B1 U$$2099/B2 VGND VGND VPWR VPWR U$$2070/A
+ sky130_fd_sc_hd__a22o_1
XU$$1335 U$$2842/A1 U$$1237/X U$$2842/B1 U$$1337/B2 VGND VGND VPWR VPWR U$$1336/A
+ sky130_fd_sc_hd__a22o_1
XU$$1346 U$$1346/A input11/X VGND VGND VPWR VPWR U$$1346/X sky130_fd_sc_hd__xor2_1
XFILLER_206_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1357 U$$946/A1 U$$1361/A2 U$$811/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1358/A sky130_fd_sc_hd__a22o_1
XFILLER_149_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1368 U$$1368/A input11/X VGND VGND VPWR VPWR U$$1368/X sky130_fd_sc_hd__xor2_1
XFILLER_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1379 U$$1379/A U$$1405/B VGND VGND VPWR VPWR U$$1379/X sky130_fd_sc_hd__xor2_1
XFILLER_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_209_ _314_/CLK _209_/D VGND VGND VPWR VPWR _209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1140 final_adder.U$$138/A final_adder.U$$847/X VGND VGND VPWR VPWR
+ output275/A sky130_fd_sc_hd__xor2_1
XFILLER_172_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1151 final_adder.U$$1151/A final_adder.U$$899/X VGND VGND VPWR VPWR
+ output287/A sky130_fd_sc_hd__xor2_2
XFILLER_156_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_51_1 dadda_fa_2_51_1/A dadda_fa_2_51_1/B dadda_fa_2_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_0/CIN dadda_fa_3_51_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_22_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_44_0 U$$2356/X U$$2489/X U$$2622/X VGND VGND VPWR VPWR dadda_fa_3_45_0/B
+ dadda_fa_3_44_2/B sky130_fd_sc_hd__fa_1
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$20 _316_/Q _188_/Q VGND VGND VPWR VPWR final_adder.U$$235/A2 final_adder.U$$234/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$31 _327_/Q _199_/Q VGND VGND VPWR VPWR final_adder.U$$225/B1 final_adder.U$$224/B
+ sky130_fd_sc_hd__ha_1
XU$$3260 U$$3260/A U$$3264/B VGND VGND VPWR VPWR U$$3260/X sky130_fd_sc_hd__xor2_1
XU$$3271 U$$3545/A1 U$$3277/A2 U$$3684/A1 U$$3277/B2 VGND VGND VPWR VPWR U$$3272/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$42 _338_/Q _210_/Q VGND VGND VPWR VPWR final_adder.U$$983/B1 final_adder.U$$212/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$53 _349_/Q _221_/Q VGND VGND VPWR VPWR final_adder.U$$203/B1 final_adder.U$$202/B
+ sky130_fd_sc_hd__ha_1
XU$$3282 U$$3282/A U$$3286/B VGND VGND VPWR VPWR U$$3282/X sky130_fd_sc_hd__xor2_1
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$64 _360_/Q _232_/Q VGND VGND VPWR VPWR final_adder.U$$961/B1 final_adder.U$$190/A
+ sky130_fd_sc_hd__ha_1
XFILLER_179_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$75 _371_/Q _243_/Q VGND VGND VPWR VPWR final_adder.U$$181/B1 final_adder.U$$180/B
+ sky130_fd_sc_hd__ha_2
XU$$3293 U$$3291/B input42/X input43/X U$$3288/Y VGND VGND VPWR VPWR U$$3293/X sky130_fd_sc_hd__a22o_4
XFILLER_59_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2570 U$$2842/B1 U$$2576/A2 U$$2709/A1 U$$2576/B2 VGND VGND VPWR VPWR U$$2571/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$86 _382_/Q _254_/Q VGND VGND VPWR VPWR final_adder.U$$939/B1 final_adder.U$$168/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$97 _393_/Q _265_/Q VGND VGND VPWR VPWR final_adder.U$$159/B1 final_adder.U$$158/B
+ sky130_fd_sc_hd__ha_1
XU$$2581 U$$2581/A U$$2602/A VGND VGND VPWR VPWR U$$2581/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2592 U$$3414/A1 U$$2600/A2 U$$3414/B1 U$$2600/B2 VGND VGND VPWR VPWR U$$2593/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1880 U$$1880/A U$$1880/B VGND VGND VPWR VPWR U$$1880/X sky130_fd_sc_hd__xor2_1
XFILLER_107_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_419 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1891 U$$2165/A1 U$$1915/A2 U$$660/A1 U$$1915/B2 VGND VGND VPWR VPWR U$$1892/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_786 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_73_2 dadda_fa_4_73_2/A dadda_fa_4_73_2/B dadda_fa_4_73_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_74_0/CIN dadda_fa_5_73_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_89_2 U$$2579/X U$$2712/X U$$2845/X VGND VGND VPWR VPWR dadda_fa_2_90_4/B
+ dadda_fa_2_89_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_66_1 dadda_fa_4_66_1/A dadda_fa_4_66_1/B dadda_fa_4_66_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/B dadda_fa_5_66_1/B sky130_fd_sc_hd__fa_1
XTAP_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_43_0 dadda_fa_7_43_0/A dadda_fa_7_43_0/B dadda_fa_7_43_0/CIN VGND VGND
+ VPWR VPWR _340_/D _211_/D sky130_fd_sc_hd__fa_2
XFILLER_77_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_59_0 dadda_fa_4_59_0/A dadda_fa_4_59_0/B dadda_fa_4_59_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/A dadda_fa_5_59_1/A sky130_fd_sc_hd__fa_1
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$510 final_adder.U$$518/B final_adder.U$$510/B VGND VGND VPWR VPWR
+ final_adder.U$$630/B sky130_fd_sc_hd__and2_1
XTAP_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$521 final_adder.U$$520/B final_adder.U$$405/X final_adder.U$$397/X
+ VGND VGND VPWR VPWR final_adder.U$$521/X sky130_fd_sc_hd__a21o_1
XTAP_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$532 final_adder.U$$540/B final_adder.U$$532/B VGND VGND VPWR VPWR
+ final_adder.U$$652/B sky130_fd_sc_hd__and2_1
XTAP_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$543 final_adder.U$$542/B final_adder.U$$427/X final_adder.U$$419/X
+ VGND VGND VPWR VPWR final_adder.U$$543/X sky130_fd_sc_hd__a21o_1
XTAP_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$554 final_adder.U$$562/B final_adder.U$$554/B VGND VGND VPWR VPWR
+ final_adder.U$$674/B sky130_fd_sc_hd__and2_1
XTAP_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$565 final_adder.U$$564/B final_adder.U$$449/X final_adder.U$$441/X
+ VGND VGND VPWR VPWR final_adder.U$$565/X sky130_fd_sc_hd__a21o_1
XTAP_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$404 U$$676/B1 U$$278/X U$$678/B1 U$$279/X VGND VGND VPWR VPWR U$$405/A sky130_fd_sc_hd__a22o_1
XFILLER_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$576 final_adder.U$$584/B final_adder.U$$576/B VGND VGND VPWR VPWR
+ final_adder.U$$696/B sky130_fd_sc_hd__and2_1
XTAP_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$415 U$$413/Y U$$412/A U$$411/A U$$414/X U$$411/Y VGND VGND VPWR VPWR U$$415/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater780 U$$2828/B2 VGND VGND VPWR VPWR U$$2874/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$587 final_adder.U$$586/B final_adder.U$$471/X final_adder.U$$463/X
+ VGND VGND VPWR VPWR final_adder.U$$587/X sky130_fd_sc_hd__a21o_1
XU$$426 U$$426/A U$$436/B VGND VGND VPWR VPWR U$$426/X sky130_fd_sc_hd__xor2_1
XTAP_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater791 U$$2600/B2 VGND VGND VPWR VPWR U$$2596/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_57_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$598 final_adder.U$$606/B final_adder.U$$598/B VGND VGND VPWR VPWR
+ final_adder.U$$718/B sky130_fd_sc_hd__and2_1
XU$$437 U$$846/B1 U$$437/A2 U$$850/A1 U$$437/B2 VGND VGND VPWR VPWR U$$438/A sky130_fd_sc_hd__a22o_1
XTAP_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$448 U$$448/A U$$474/B VGND VGND VPWR VPWR U$$448/X sky130_fd_sc_hd__xor2_1
XFILLER_72_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$459 U$$594/B1 U$$491/A2 U$$461/A1 U$$491/B2 VGND VGND VPWR VPWR U$$460/A sky130_fd_sc_hd__a22o_1
XFILLER_44_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4423_1788 VGND VGND VPWR VPWR U$$4423_1788/HI U$$4423/B sky130_fd_sc_hd__conb_1
XFILLER_139_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1304 U$$3425/A VGND VGND VPWR VPWR U$$3349/B sky130_fd_sc_hd__buf_8
Xrepeater1315 U$$3244/B VGND VGND VPWR VPWR U$$3228/B sky130_fd_sc_hd__buf_6
Xrepeater1326 U$$3133/B VGND VGND VPWR VPWR U$$3150/A sky130_fd_sc_hd__buf_8
XFILLER_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1337 U$$3008/B VGND VGND VPWR VPWR U$$3013/A sky130_fd_sc_hd__buf_6
XFILLER_176_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1348 input36/X VGND VGND VPWR VPWR U$$2845/B sky130_fd_sc_hd__buf_6
XFILLER_5_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1359 U$$2658/B VGND VGND VPWR VPWR U$$2624/B sky130_fd_sc_hd__clkbuf_8
XFILLER_84_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_842 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_61_0 dadda_fa_3_61_0/A dadda_fa_3_61_0/B dadda_fa_3_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_0/B dadda_fa_4_61_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_77_0 U$$958/Y U$$1092/X U$$1225/X VGND VGND VPWR VPWR dadda_fa_1_78_8/CIN
+ dadda_fa_2_77_0/A sky130_fd_sc_hd__fa_1
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_ha_4_8_0 U$$23/X U$$156/X VGND VGND VPWR VPWR dadda_fa_5_9_1/B dadda_ha_4_8_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$960 input6/X VGND VGND VPWR VPWR U$$962/B sky130_fd_sc_hd__inv_1
XU$$971 U$$12/A1 U$$979/A2 U$$14/A1 U$$979/B2 VGND VGND VPWR VPWR U$$972/A sky130_fd_sc_hd__a22o_1
XU$$1110 U$$2069/A1 U$$1138/A2 U$$2206/B1 U$$1138/B2 VGND VGND VPWR VPWR U$$1111/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1121 U$$1121/A U$$1137/B VGND VGND VPWR VPWR U$$1121/X sky130_fd_sc_hd__xor2_1
XU$$982 U$$982/A U$$996/B VGND VGND VPWR VPWR U$$982/X sky130_fd_sc_hd__xor2_1
XFILLER_62_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1132 U$$719/B1 U$$1136/A2 U$$721/B1 U$$1136/B2 VGND VGND VPWR VPWR U$$1133/A sky130_fd_sc_hd__a22o_1
XFILLER_204_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$993 U$$993/A1 U$$993/A2 U$$993/B1 U$$993/B2 VGND VGND VPWR VPWR U$$994/A sky130_fd_sc_hd__a22o_1
XFILLER_44_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_662 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1143 U$$1143/A U$$1187/B VGND VGND VPWR VPWR U$$1143/X sky130_fd_sc_hd__xor2_1
XFILLER_210_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1154 U$$58/A1 U$$1162/A2 U$$60/A1 U$$1162/B2 VGND VGND VPWR VPWR U$$1155/A sky130_fd_sc_hd__a22o_1
XFILLER_188_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1165 U$$1165/A U$$1187/B VGND VGND VPWR VPWR U$$1165/X sky130_fd_sc_hd__xor2_1
XFILLER_203_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1176 U$$902/A1 U$$1222/A2 U$$4055/A1 U$$1222/B2 VGND VGND VPWR VPWR U$$1177/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1187 U$$1187/A U$$1187/B VGND VGND VPWR VPWR U$$1187/X sky130_fd_sc_hd__xor2_1
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1198 U$$2842/A1 U$$1204/A2 U$$2842/B1 U$$1204/B2 VGND VGND VPWR VPWR U$$1199/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_83_1 dadda_fa_5_83_1/A dadda_fa_5_83_1/B dadda_fa_5_83_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_84_0/B dadda_fa_7_83_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_2_99_1 U$$2865/X U$$2998/X U$$3131/X VGND VGND VPWR VPWR dadda_fa_3_100_1/B
+ dadda_fa_3_99_3/A sky130_fd_sc_hd__fa_1
XFILLER_172_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_76_0 dadda_fa_5_76_0/A dadda_fa_5_76_0/B dadda_fa_5_76_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_77_0/A dadda_fa_6_76_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_75_8 dadda_fa_1_75_8/A dadda_fa_1_75_8/B dadda_fa_1_75_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_76_3/A dadda_fa_3_75_0/A sky130_fd_sc_hd__fa_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_68_7 dadda_fa_1_68_7/A dadda_fa_1_68_7/B dadda_fa_1_68_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_2/CIN dadda_fa_2_68_5/CIN sky130_fd_sc_hd__fa_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3090 input92/X U$$3118/A2 U$$4049/B1 U$$3118/B2 VGND VGND VPWR VPWR U$$3091/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_399 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_94_0 dadda_fa_1_94_0/A U$$2190/X U$$2323/X VGND VGND VPWR VPWR dadda_fa_2_95_5/B
+ dadda_fa_2_94_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_2_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$340 final_adder.U$$342/B final_adder.U$$340/B VGND VGND VPWR VPWR
+ final_adder.U$$466/B sky130_fd_sc_hd__and2_1
XTAP_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$351 final_adder.U$$350/B final_adder.U$$225/X final_adder.U$$223/X
+ VGND VGND VPWR VPWR final_adder.U$$351/X sky130_fd_sc_hd__a21o_1
XTAP_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_106_0 dadda_fa_6_106_0/A dadda_fa_6_106_0/B dadda_fa_6_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_107_0/B dadda_fa_7_106_0/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$362 final_adder.U$$364/B final_adder.U$$362/B VGND VGND VPWR VPWR
+ final_adder.U$$488/B sky130_fd_sc_hd__and2_1
XTAP_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$201 U$$64/A1 U$$259/A2 U$$66/A1 U$$259/B2 VGND VGND VPWR VPWR U$$202/A sky130_fd_sc_hd__a22o_1
XTAP_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$373 final_adder.U$$372/B final_adder.U$$247/X final_adder.U$$245/X
+ VGND VGND VPWR VPWR final_adder.U$$373/X sky130_fd_sc_hd__a21o_1
XTAP_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$212 U$$212/A U$$212/B VGND VGND VPWR VPWR U$$212/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$384 final_adder.U$$388/B final_adder.U$$384/B VGND VGND VPWR VPWR
+ final_adder.U$$508/B sky130_fd_sc_hd__and2_1
XTAP_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$223 U$$86/A1 U$$263/A2 U$$88/A1 U$$231/B2 VGND VGND VPWR VPWR U$$224/A sky130_fd_sc_hd__a22o_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$395 final_adder.U$$394/B final_adder.U$$273/X final_adder.U$$269/X
+ VGND VGND VPWR VPWR final_adder.U$$395/X sky130_fd_sc_hd__a21o_1
XTAP_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$234 U$$234/A U$$244/B VGND VGND VPWR VPWR U$$234/X sky130_fd_sc_hd__xor2_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$245 U$$654/B1 U$$257/A2 U$$521/A1 U$$257/B2 VGND VGND VPWR VPWR U$$246/A sky130_fd_sc_hd__a22o_1
XTAP_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$256 U$$256/A U$$260/B VGND VGND VPWR VPWR U$$256/X sky130_fd_sc_hd__xor2_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_26_3 dadda_fa_3_26_3/A dadda_fa_3_26_3/B dadda_fa_3_26_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_27_1/B dadda_fa_4_26_2/CIN sky130_fd_sc_hd__fa_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$267 U$$676/B1 U$$141/X U$$678/B1 U$$142/X VGND VGND VPWR VPWR U$$268/A sky130_fd_sc_hd__a22o_1
XFILLER_72_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$278 U$$276/Y U$$275/A U$$274/A U$$277/X U$$274/Y VGND VGND VPWR VPWR U$$278/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$289 U$$289/A U$$317/B VGND VGND VPWR VPWR U$$289/X sky130_fd_sc_hd__xor2_1
XFILLER_26_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_1209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_93_0 dadda_fa_6_93_0/A dadda_fa_6_93_0/B dadda_fa_6_93_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_94_0/B dadda_fa_7_93_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_139_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$6 U$$6/A1 U$$8/A2 U$$8/A1 U$$8/B2 VGND VGND VPWR VPWR U$$7/A sky130_fd_sc_hd__a22o_1
XFILLER_126_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1101 U$$3296/B1 VGND VGND VPWR VPWR U$$2202/A1 sky130_fd_sc_hd__buf_6
XFILLER_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1112 U$$4019/A1 VGND VGND VPWR VPWR U$$3880/B1 sky130_fd_sc_hd__buf_8
Xoutput309 output309/A VGND VGND VPWR VPWR o[31] sky130_fd_sc_hd__buf_2
Xrepeater1123 U$$4013/B1 VGND VGND VPWR VPWR U$$179/A1 sky130_fd_sc_hd__buf_4
XFILLER_126_455 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1134 U$$4424/A1 VGND VGND VPWR VPWR U$$4011/B1 sky130_fd_sc_hd__buf_6
Xrepeater1145 input71/X VGND VGND VPWR VPWR U$$4422/A1 sky130_fd_sc_hd__buf_12
XFILLER_126_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1156 U$$998/B VGND VGND VPWR VPWR U$$980/B sky130_fd_sc_hd__buf_6
Xrepeater1167 U$$4144/A1 VGND VGND VPWR VPWR U$$3183/B1 sky130_fd_sc_hd__buf_6
Xrepeater1178 input68/X VGND VGND VPWR VPWR U$$32/A1 sky130_fd_sc_hd__buf_4
XFILLER_206_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1189 U$$850/A1 VGND VGND VPWR VPWR U$$987/A1 sky130_fd_sc_hd__buf_6
XFILLER_171_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$790 U$$790/A U$$821/A VGND VGND VPWR VPWR U$$790/X sky130_fd_sc_hd__xor2_1
XFILLER_16_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1099 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_411 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_80_6 U$$3492/X U$$3625/X U$$3758/X VGND VGND VPWR VPWR dadda_fa_2_81_2/CIN
+ dadda_fa_2_80_5/B sky130_fd_sc_hd__fa_1
Xrepeater1690 U$$3245/A1 VGND VGND VPWR VPWR U$$2834/A1 sky130_fd_sc_hd__buf_6
XFILLER_104_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_73_5 U$$3877/X U$$4010/X U$$4143/X VGND VGND VPWR VPWR dadda_fa_2_74_2/A
+ dadda_fa_2_73_5/A sky130_fd_sc_hd__fa_1
XFILLER_58_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_66_4 U$$4129/X U$$4262/X U$$4395/X VGND VGND VPWR VPWR dadda_fa_2_67_1/CIN
+ dadda_fa_2_66_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_59_3 U$$2785/X U$$2918/X U$$3051/X VGND VGND VPWR VPWR dadda_fa_2_60_1/B
+ dadda_fa_2_59_4/B sky130_fd_sc_hd__fa_1
XFILLER_100_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_36_2 dadda_fa_4_36_2/A dadda_fa_4_36_2/B dadda_fa_4_36_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_37_0/CIN dadda_fa_5_36_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_29_1 dadda_fa_4_29_1/A dadda_fa_4_29_1/B dadda_fa_4_29_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/B dadda_fa_5_29_1/B sky130_fd_sc_hd__fa_1
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_469 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_190_ _326_/CLK _190_/D VGND VGND VPWR VPWR _190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_528 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_0_62_5 U$$2126/X U$$2259/X VGND VGND VPWR VPWR dadda_fa_1_63_7/A dadda_fa_2_62_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_68_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$4505 U$$4505/A U$$4505/B VGND VGND VPWR VPWR U$$4505/X sky130_fd_sc_hd__xor2_1
XU$$4516 U$$4516/A1 U$$4388/X U$$4516/B1 U$$4389/X VGND VGND VPWR VPWR U$$4517/A sky130_fd_sc_hd__a22o_1
XTAP_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_61_3 U$$1326/X U$$1459/X U$$1592/X VGND VGND VPWR VPWR dadda_fa_1_62_6/CIN
+ dadda_fa_1_61_8/CIN sky130_fd_sc_hd__fa_1
XTAP_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3804 U$$3804/A U$$3826/B VGND VGND VPWR VPWR U$$3804/X sky130_fd_sc_hd__xor2_1
XU$$19 U$$19/A U$$43/B VGND VGND VPWR VPWR U$$19/X sky130_fd_sc_hd__xor2_1
XFILLER_18_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3815 U$$4361/B1 U$$3819/A2 U$$4228/A1 U$$3819/B2 VGND VGND VPWR VPWR U$$3816/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3826 U$$3826/A U$$3826/B VGND VGND VPWR VPWR U$$3826/X sky130_fd_sc_hd__xor2_1
XFILLER_131_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3837 input52/X VGND VGND VPWR VPWR U$$3839/B sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$170 final_adder.U$$170/A final_adder.U$$170/B VGND VGND VPWR VPWR
+ final_adder.U$$298/B sky130_fd_sc_hd__and2_1
XTAP_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$181 final_adder.U$$180/B final_adder.U$$951/B1 final_adder.U$$181/B1
+ VGND VGND VPWR VPWR final_adder.U$$181/X sky130_fd_sc_hd__a21o_1
XTAP_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_31_1 dadda_fa_3_31_1/A dadda_fa_3_31_1/B dadda_fa_3_31_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_0/CIN dadda_fa_4_31_2/A sky130_fd_sc_hd__fa_1
XU$$3848 input87/X U$$3878/A2 input98/X U$$3878/B2 VGND VGND VPWR VPWR U$$3849/A sky130_fd_sc_hd__a22o_1
XTAP_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3859 U$$3859/A U$$3875/B VGND VGND VPWR VPWR U$$3859/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$192 final_adder.U$$192/A final_adder.U$$192/B VGND VGND VPWR VPWR
+ final_adder.U$$320/B sky130_fd_sc_hd__and2_1
XFILLER_166_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_24_0 U$$720/X U$$853/X U$$986/X VGND VGND VPWR VPWR dadda_fa_4_25_0/B
+ dadda_fa_4_24_1/CIN sky130_fd_sc_hd__fa_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_388_ _421_/CLK _388_/D VGND VGND VPWR VPWR _388_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1102 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_90_5 dadda_fa_2_90_5/A dadda_fa_2_90_5/B dadda_fa_2_90_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_91_2/A dadda_fa_4_90_0/A sky130_fd_sc_hd__fa_2
XFILLER_138_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_403 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_83_4 dadda_fa_2_83_4/A dadda_fa_2_83_4/B dadda_fa_2_83_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_1/CIN dadda_fa_3_83_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_76_3 dadda_fa_2_76_3/A dadda_fa_2_76_3/B dadda_fa_2_76_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/B dadda_fa_3_76_3/B sky130_fd_sc_hd__fa_1
XFILLER_68_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_69_2 dadda_fa_2_69_2/A dadda_fa_2_69_2/B dadda_fa_2_69_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/A dadda_fa_3_69_3/A sky130_fd_sc_hd__fa_2
XFILLER_96_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_46_1 dadda_fa_5_46_1/A dadda_fa_5_46_1/B dadda_fa_5_46_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_47_0/B dadda_fa_7_46_0/A sky130_fd_sc_hd__fa_1
XFILLER_56_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_39_0 dadda_fa_5_39_0/A dadda_fa_5_39_0/B dadda_fa_5_39_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_40_0/A dadda_fa_6_39_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_3_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_832 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_120_1 dadda_fa_5_120_1/A dadda_fa_5_120_1/B dadda_ha_4_120_1/SUM VGND
+ VGND VPWR VPWR dadda_fa_6_121_0/B dadda_fa_7_120_0/A sky130_fd_sc_hd__fa_1
XFILLER_164_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_113_0 dadda_fa_5_113_0/A dadda_fa_5_113_0/B dadda_fa_5_113_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_114_0/A dadda_fa_6_113_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_71_2 U$$2942/X U$$3075/X U$$3208/X VGND VGND VPWR VPWR dadda_fa_2_72_1/A
+ dadda_fa_2_71_4/A sky130_fd_sc_hd__fa_1
XFILLER_154_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_1 U$$2928/X U$$3061/X U$$3194/X VGND VGND VPWR VPWR dadda_fa_2_65_0/CIN
+ dadda_fa_2_64_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_41_0 dadda_fa_4_41_0/A dadda_fa_4_41_0/B dadda_fa_4_41_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/A dadda_fa_5_41_1/A sky130_fd_sc_hd__fa_1
XFILLER_115_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_57_0 U$$1185/X U$$1318/X U$$1451/X VGND VGND VPWR VPWR dadda_fa_2_58_0/B
+ dadda_fa_2_57_3/B sky130_fd_sc_hd__fa_1
XFILLER_41_1263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1709 U$$1709/A U$$1721/B VGND VGND VPWR VPWR U$$1709/X sky130_fd_sc_hd__xor2_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_311_ _337_/CLK _311_/D VGND VGND VPWR VPWR _311_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_242_ _246_/CLK _242_/D VGND VGND VPWR VPWR _242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_173_ _304_/CLK _173_/D VGND VGND VPWR VPWR _173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput19 a[26] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_196_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_93_3 dadda_fa_3_93_3/A dadda_fa_3_93_3/B dadda_fa_3_93_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_94_1/B dadda_fa_4_93_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_86_2 dadda_fa_3_86_2/A dadda_fa_3_86_2/B dadda_fa_3_86_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_1/A dadda_fa_4_86_2/B sky130_fd_sc_hd__fa_1
XFILLER_184_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_79_1 dadda_fa_3_79_1/A dadda_fa_3_79_1/B dadda_fa_3_79_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_0/CIN dadda_fa_4_79_2/A sky130_fd_sc_hd__fa_1
XFILLER_69_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_56_0 dadda_fa_6_56_0/A dadda_fa_6_56_0/B dadda_fa_6_56_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_57_0/B dadda_fa_7_56_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_151_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1005 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater609 U$$175/A2 VGND VGND VPWR VPWR U$$165/A2 sky130_fd_sc_hd__buf_2
XFILLER_81_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4302 U$$4302/A U$$4384/A VGND VGND VPWR VPWR U$$4302/X sky130_fd_sc_hd__xor2_1
XU$$4313 input86/X U$$4361/A2 input88/X U$$4361/B2 VGND VGND VPWR VPWR U$$4314/A sky130_fd_sc_hd__a22o_1
XFILLER_42_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_364 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4324 U$$4324/A U$$4330/B VGND VGND VPWR VPWR U$$4324/X sky130_fd_sc_hd__xor2_1
XU$$4335 input99/X U$$4349/A2 U$$4335/B1 U$$4349/B2 VGND VGND VPWR VPWR U$$4336/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4346 U$$4346/A U$$4366/B VGND VGND VPWR VPWR U$$4346/X sky130_fd_sc_hd__xor2_1
XU$$3601 U$$3601/A U$$3637/B VGND VGND VPWR VPWR U$$3601/X sky130_fd_sc_hd__xor2_1
XFILLER_203_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4357 input111/X U$$4373/A2 U$$4496/A1 U$$4373/B2 VGND VGND VPWR VPWR U$$4358/A
+ sky130_fd_sc_hd__a22o_1
XU$$3612 U$$3884/B1 U$$3612/A2 U$$3612/B1 U$$3612/B2 VGND VGND VPWR VPWR U$$3613/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_115_2 dadda_fa_4_115_2/A dadda_fa_4_115_2/B dadda_fa_4_115_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_116_0/CIN dadda_fa_5_115_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3623 U$$3623/A U$$3623/B VGND VGND VPWR VPWR U$$3623/X sky130_fd_sc_hd__xor2_1
XU$$4368 U$$4368/A U$$4370/B VGND VGND VPWR VPWR U$$4368/X sky130_fd_sc_hd__xor2_1
XU$$3634 U$$4043/B1 U$$3636/A2 U$$3908/B1 U$$3636/B2 VGND VGND VPWR VPWR U$$3635/A
+ sky130_fd_sc_hd__a22o_1
XU$$4379 U$$4379/A1 U$$4251/X U$$4516/B1 U$$4252/X VGND VGND VPWR VPWR U$$4380/A sky130_fd_sc_hd__a22o_1
XFILLER_18_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3645 U$$3645/A U$$3697/B VGND VGND VPWR VPWR U$$3645/X sky130_fd_sc_hd__xor2_1
XU$$2900 U$$2900/A U$$2920/B VGND VGND VPWR VPWR U$$2900/X sky130_fd_sc_hd__xor2_1
XU$$2911 U$$32/B1 U$$2919/A2 U$$4146/A1 U$$2919/B2 VGND VGND VPWR VPWR U$$2912/A sky130_fd_sc_hd__a22o_1
XU$$3656 U$$4476/B1 U$$3660/A2 U$$4343/A1 U$$3660/B2 VGND VGND VPWR VPWR U$$3657/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_108_1 dadda_fa_4_108_1/A dadda_fa_4_108_1/B dadda_fa_4_108_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/B dadda_fa_5_108_1/B sky130_fd_sc_hd__fa_1
XFILLER_19_987 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2922 U$$2922/A U$$2922/B VGND VGND VPWR VPWR U$$2922/X sky130_fd_sc_hd__xor2_1
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3667 U$$3667/A U$$3683/B VGND VGND VPWR VPWR U$$3667/X sky130_fd_sc_hd__xor2_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3678 U$$388/B1 U$$3680/A2 U$$3817/A1 U$$3680/B2 VGND VGND VPWR VPWR U$$3679/A
+ sky130_fd_sc_hd__a22o_1
XU$$2933 U$$4440/A1 U$$2977/A2 U$$4440/B1 U$$2979/B2 VGND VGND VPWR VPWR U$$2934/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3689 U$$3689/A U$$3698/A VGND VGND VPWR VPWR U$$3689/X sky130_fd_sc_hd__xor2_1
XFILLER_34_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2944 U$$2944/A U$$2968/B VGND VGND VPWR VPWR U$$2944/X sky130_fd_sc_hd__xor2_1
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2955 U$$2955/A1 U$$2985/A2 U$$2957/A1 U$$2985/B2 VGND VGND VPWR VPWR U$$2956/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_946 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2966 U$$2966/A U$$2978/B VGND VGND VPWR VPWR U$$2966/X sky130_fd_sc_hd__xor2_1
XU$$2977 U$$3114/A1 U$$2977/A2 U$$3116/A1 U$$2882/X VGND VGND VPWR VPWR U$$2978/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 U$$2052/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2988 U$$2988/A U$$2996/B VGND VGND VPWR VPWR U$$2988/X sky130_fd_sc_hd__xor2_1
XANTENNA_271 U$$1746/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2999 U$$122/A1 U$$3011/A2 U$$3547/B1 U$$3011/B2 VGND VGND VPWR VPWR U$$3000/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_158_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_859 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$691_1841 VGND VGND VPWR VPWR U$$691_1841/HI U$$691/A1 sky130_fd_sc_hd__conb_1
XFILLER_127_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1071 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_81_1 dadda_fa_2_81_1/A dadda_fa_2_81_1/B dadda_fa_2_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_0/CIN dadda_fa_3_81_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_64_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_74_0 dadda_fa_2_74_0/A dadda_fa_2_74_0/B dadda_fa_2_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_0/B dadda_fa_3_74_2/B sky130_fd_sc_hd__fa_1
XFILLER_130_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$917 final_adder.U$$146/A final_adder.U$$855/X final_adder.U$$917/B1
+ VGND VGND VPWR VPWR final_adder.U$$917/X sky130_fd_sc_hd__a21o_1
XFILLER_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$939 final_adder.U$$168/A final_adder.U$$877/X final_adder.U$$939/B1
+ VGND VGND VPWR VPWR final_adder.U$$939/X sky130_fd_sc_hd__a21o_1
XFILLER_56_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_50_7 U$$2900/X U$$3033/X U$$3166/X VGND VGND VPWR VPWR dadda_fa_2_51_2/CIN
+ dadda_fa_2_50_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_113_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_740 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_607 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_787 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_96_1 dadda_fa_4_96_1/A dadda_fa_4_96_1/B dadda_fa_4_96_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/B dadda_fa_5_96_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_7_73_0 dadda_fa_7_73_0/A dadda_fa_7_73_0/B dadda_fa_7_73_0/CIN VGND VGND
+ VPWR VPWR _370_/D _241_/D sky130_fd_sc_hd__fa_1
Xdadda_fa_4_89_0 dadda_fa_4_89_0/A dadda_fa_4_89_0/B dadda_fa_4_89_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/A dadda_fa_5_89_1/A sky130_fd_sc_hd__fa_1
XFILLER_69_1152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2207 U$$2207/A U$$2227/B VGND VGND VPWR VPWR U$$2207/X sky130_fd_sc_hd__xor2_1
XU$$2218 U$$2492/A1 U$$2272/A2 U$$2220/A1 U$$2272/B2 VGND VGND VPWR VPWR U$$2219/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2229 U$$2229/A U$$2253/B VGND VGND VPWR VPWR U$$2229/X sky130_fd_sc_hd__xor2_1
XU$$1506 U$$1506/A VGND VGND VPWR VPWR U$$1506/Y sky130_fd_sc_hd__inv_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1517 U$$2063/B1 U$$1545/A2 U$$2065/B1 U$$1545/B2 VGND VGND VPWR VPWR U$$1518/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1528 U$$1528/A U$$1546/B VGND VGND VPWR VPWR U$$1528/X sky130_fd_sc_hd__xor2_1
XFILLER_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1539 U$$854/A1 U$$1575/A2 U$$854/B1 U$$1575/B2 VGND VGND VPWR VPWR U$$1540/A sky130_fd_sc_hd__a22o_1
XFILLER_203_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_910 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_225_ _355_/CLK _225_/D VGND VGND VPWR VPWR _225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_91_0 dadda_fa_3_91_0/A dadda_fa_3_91_0/B dadda_fa_3_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_0/B dadda_fa_4_91_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_137_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater406 U$$689/X VGND VGND VPWR VPWR U$$805/A2 sky130_fd_sc_hd__buf_6
XFILLER_66_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater417 U$$4251/X VGND VGND VPWR VPWR U$$4381/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater428 U$$491/A2 VGND VGND VPWR VPWR U$$483/A2 sky130_fd_sc_hd__buf_6
XU$$4110 U$$4110/A VGND VGND VPWR VPWR U$$4110/Y sky130_fd_sc_hd__inv_1
Xdadda_fa_2_53_5 dadda_fa_2_53_5/A dadda_fa_2_53_5/B dadda_fa_2_53_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_54_2/A dadda_fa_4_53_0/A sky130_fd_sc_hd__fa_1
Xrepeater439 U$$94/A2 VGND VGND VPWR VPWR U$$98/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_4_120_0 dadda_fa_4_120_0/A U$$3971/X U$$4104/X VGND VGND VPWR VPWR dadda_fa_5_121_1/A
+ dadda_fa_5_120_1/B sky130_fd_sc_hd__fa_1
XFILLER_120_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4121 U$$4121/A U$$4145/B VGND VGND VPWR VPWR U$$4121/X sky130_fd_sc_hd__xor2_1
XFILLER_65_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4132 U$$4406/A1 U$$4164/A2 U$$4408/A1 U$$4164/B2 VGND VGND VPWR VPWR U$$4133/A
+ sky130_fd_sc_hd__a22o_1
XU$$4143 U$$4143/A U$$4145/B VGND VGND VPWR VPWR U$$4143/X sky130_fd_sc_hd__xor2_1
XU$$4154 input74/X U$$4188/A2 input75/X U$$4188/B2 VGND VGND VPWR VPWR U$$4155/A sky130_fd_sc_hd__a22o_1
XU$$3420 input123/X U$$3422/A2 input124/X U$$3422/B2 VGND VGND VPWR VPWR U$$3421/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_46_4 dadda_fa_2_46_4/A dadda_fa_2_46_4/B dadda_fa_2_46_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_1/CIN dadda_fa_3_46_3/CIN sky130_fd_sc_hd__fa_1
XU$$4165 U$$4165/A U$$4165/B VGND VGND VPWR VPWR U$$4165/X sky130_fd_sc_hd__xor2_1
XU$$3431 U$$3431/A1 U$$3453/A2 input65/X U$$3453/B2 VGND VGND VPWR VPWR U$$3432/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4176 U$$4176/A1 U$$4176/A2 U$$4176/B1 U$$4176/B2 VGND VGND VPWR VPWR U$$4177/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3442 U$$3442/A U$$3528/B VGND VGND VPWR VPWR U$$3442/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4187 U$$4187/A U$$4189/B VGND VGND VPWR VPWR U$$4187/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4198 U$$4333/B1 U$$4210/A2 input100/X U$$4210/B2 VGND VGND VPWR VPWR U$$4199/A
+ sky130_fd_sc_hd__a22o_1
XU$$3453 U$$3453/A1 U$$3453/A2 U$$3727/B1 U$$3453/B2 VGND VGND VPWR VPWR U$$3454/A
+ sky130_fd_sc_hd__a22o_1
XU$$3464 U$$3464/A U$$3504/B VGND VGND VPWR VPWR U$$3464/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_39_3 U$$2346/X U$$2479/X U$$2612/X VGND VGND VPWR VPWR dadda_fa_3_40_1/B
+ dadda_fa_3_39_3/B sky130_fd_sc_hd__fa_1
XU$$2730 U$$2730/A U$$2736/B VGND VGND VPWR VPWR U$$2730/X sky130_fd_sc_hd__xor2_1
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3475 U$$3884/B1 U$$3479/A2 U$$4162/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3476/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2741 input35/X VGND VGND VPWR VPWR U$$2743/B sky130_fd_sc_hd__inv_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3486 U$$3486/A U$$3490/B VGND VGND VPWR VPWR U$$3486/X sky130_fd_sc_hd__xor2_1
XU$$2752 U$$3026/A1 U$$2796/A2 U$$3028/A1 U$$2796/B2 VGND VGND VPWR VPWR U$$2753/A
+ sky130_fd_sc_hd__a22o_1
XU$$3497 U$$4043/B1 U$$3503/A2 U$$3908/B1 U$$3503/B2 VGND VGND VPWR VPWR U$$3498/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2763 U$$2763/A U$$2783/B VGND VGND VPWR VPWR U$$2763/X sky130_fd_sc_hd__xor2_1
XFILLER_179_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2774 U$$32/B1 U$$2868/A2 U$$4146/A1 U$$2868/B2 VGND VGND VPWR VPWR U$$2775/A sky130_fd_sc_hd__a22o_1
XFILLER_34_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2785 U$$2785/A U$$2817/B VGND VGND VPWR VPWR U$$2785/X sky130_fd_sc_hd__xor2_1
XU$$2796 U$$3344/A1 U$$2796/A2 U$$3207/B1 U$$2796/B2 VGND VGND VPWR VPWR U$$2797/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1078 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_689 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4451_1802 VGND VGND VPWR VPWR U$$4451_1802/HI U$$4451/B sky130_fd_sc_hd__conb_1
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput209 c[57] VGND VGND VPWR VPWR input209/X sky130_fd_sc_hd__clkbuf_4
XTAP_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$703 final_adder.U$$702/B final_adder.U$$599/X final_adder.U$$583/X
+ VGND VGND VPWR VPWR final_adder.U$$703/X sky130_fd_sc_hd__a21o_1
XTAP_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$714 final_adder.U$$714/A final_adder.U$$714/B VGND VGND VPWR VPWR
+ final_adder.U$$794/A sky130_fd_sc_hd__and2_1
XFILLER_25_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$725 final_adder.U$$708/A final_adder.U$$621/X final_adder.U$$605/X
+ VGND VGND VPWR VPWR final_adder.U$$725/X sky130_fd_sc_hd__a21o_2
Xrepeater940 input95/X VGND VGND VPWR VPWR U$$3368/B1 sky130_fd_sc_hd__buf_6
XFILLER_112_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$747 final_adder.U$$746/B final_adder.U$$667/X final_adder.U$$635/X
+ VGND VGND VPWR VPWR final_adder.U$$747/X sky130_fd_sc_hd__a21o_1
XFILLER_68_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater951 U$$4323/B1 VGND VGND VPWR VPWR U$$78/A1 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$758 final_adder.U$$790/B final_adder.U$$758/B VGND VGND VPWR VPWR
+ final_adder.U$$758/X sky130_fd_sc_hd__and2_1
Xrepeater962 U$$896/B1 VGND VGND VPWR VPWR U$$759/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_56_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$769 final_adder.U$$768/B final_adder.U$$689/X final_adder.U$$657/X
+ VGND VGND VPWR VPWR final_adder.U$$769/X sky130_fd_sc_hd__a21o_1
XU$$608 U$$745/A1 U$$636/A2 U$$610/A1 U$$636/B2 VGND VGND VPWR VPWR U$$609/A sky130_fd_sc_hd__a22o_1
Xrepeater973 input91/X VGND VGND VPWR VPWR U$$3908/B1 sky130_fd_sc_hd__buf_4
XFILLER_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$619 U$$619/A U$$625/B VGND VGND VPWR VPWR U$$619/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater984 U$$1175/B VGND VGND VPWR VPWR U$$1139/B sky130_fd_sc_hd__buf_6
Xrepeater995 input89/X VGND VGND VPWR VPWR U$$4454/A1 sky130_fd_sc_hd__buf_4
XFILLER_17_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_409 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1508 U$$3829/A1 VGND VGND VPWR VPWR U$$952/A1 sky130_fd_sc_hd__buf_4
XFILLER_116_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1519 U$$4099/B1 VGND VGND VPWR VPWR U$$4512/A1 sky130_fd_sc_hd__buf_6
XFILLER_193_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_108_0 U$$3282/X U$$3415/X U$$3548/X VGND VGND VPWR VPWR dadda_fa_4_109_0/B
+ dadda_fa_4_108_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_919 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_56_3 dadda_fa_3_56_3/A dadda_fa_3_56_3/B dadda_fa_3_56_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_57_1/B dadda_fa_4_56_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_49_2 dadda_fa_3_49_2/A dadda_fa_3_49_2/B dadda_fa_3_49_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_1/A dadda_fa_4_49_2/B sky130_fd_sc_hd__fa_1
XFILLER_208_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2004 U$$3235/B1 U$$2022/A2 U$$2691/A1 U$$2022/B2 VGND VGND VPWR VPWR U$$2005/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2015 U$$2015/A U$$2037/B VGND VGND VPWR VPWR U$$2015/X sky130_fd_sc_hd__xor2_1
XFILLER_63_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_19_0 dadda_fa_6_19_0/A dadda_fa_6_19_0/B dadda_fa_6_19_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_20_0/B dadda_fa_7_19_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2026 U$$2026/A1 U$$2052/A2 U$$930/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2027/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2037 U$$2037/A U$$2037/B VGND VGND VPWR VPWR U$$2037/X sky130_fd_sc_hd__xor2_1
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2048 U$$4375/B1 U$$2052/A2 U$$4103/B1 U$$2052/B2 VGND VGND VPWR VPWR U$$2049/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1303 U$$70/A1 U$$1323/A2 U$$72/A1 U$$1307/B2 VGND VGND VPWR VPWR U$$1304/A sky130_fd_sc_hd__a22o_1
XU$$1314 U$$1314/A U$$1316/B VGND VGND VPWR VPWR U$$1314/X sky130_fd_sc_hd__xor2_1
XU$$2059 U$$2057/Y input24/X input22/X U$$2058/X U$$2055/Y VGND VGND VPWR VPWR U$$2059/X
+ sky130_fd_sc_hd__a32o_2
XU$$1325 U$$92/A1 U$$1337/A2 U$$94/A1 U$$1337/B2 VGND VGND VPWR VPWR U$$1326/A sky130_fd_sc_hd__a22o_1
XFILLER_15_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1336 U$$1336/A U$$1338/B VGND VGND VPWR VPWR U$$1336/X sky130_fd_sc_hd__xor2_1
XFILLER_16_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1347 U$$799/A1 U$$1367/A2 U$$2582/A1 U$$1367/B2 VGND VGND VPWR VPWR U$$1348/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1358 U$$1358/A U$$1366/B VGND VGND VPWR VPWR U$$1358/X sky130_fd_sc_hd__xor2_1
XFILLER_206_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1369 input11/X VGND VGND VPWR VPWR U$$1369/Y sky130_fd_sc_hd__inv_1
XFILLER_43_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_208_ _208_/CLK _208_/D VGND VGND VPWR VPWR _208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1130 final_adder.U$$148/A final_adder.U$$857/X VGND VGND VPWR VPWR
+ output264/A sky130_fd_sc_hd__xor2_1
XFILLER_190_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1141 final_adder.U$$138/B final_adder.U$$909/X VGND VGND VPWR VPWR
+ output276/A sky130_fd_sc_hd__xor2_1
XFILLER_128_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_51_2 dadda_fa_2_51_2/A dadda_fa_2_51_2/B dadda_fa_2_51_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/A dadda_fa_3_51_3/A sky130_fd_sc_hd__fa_1
XFILLER_22_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_44_1 U$$2755/X U$$2888/X U$$3021/X VGND VGND VPWR VPWR dadda_fa_3_45_0/CIN
+ dadda_fa_3_44_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_66_665 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$10 _306_/Q _178_/Q VGND VGND VPWR VPWR final_adder.U$$245/A2 final_adder.U$$244/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$21 _317_/Q _189_/Q VGND VGND VPWR VPWR final_adder.U$$235/B1 final_adder.U$$234/B
+ sky130_fd_sc_hd__ha_1
XU$$4481_1817 VGND VGND VPWR VPWR U$$4481_1817/HI U$$4481/B sky130_fd_sc_hd__conb_1
XU$$3250 U$$3250/A U$$3286/B VGND VGND VPWR VPWR U$$3250/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_21_0 dadda_fa_5_21_0/A dadda_fa_5_21_0/B dadda_fa_5_21_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_22_0/A dadda_fa_6_21_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_54_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$32 _328_/Q _200_/Q VGND VGND VPWR VPWR final_adder.U$$993/B1 final_adder.U$$222/A
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_2_37_0 U$$746/X U$$879/X U$$1012/X VGND VGND VPWR VPWR dadda_fa_3_38_0/B
+ dadda_fa_3_37_2/B sky130_fd_sc_hd__fa_1
XFILLER_81_635 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3261 U$$521/A1 U$$3263/A2 U$$384/B1 U$$3263/B2 VGND VGND VPWR VPWR U$$3262/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$43 _339_/Q _211_/Q VGND VGND VPWR VPWR final_adder.U$$213/B1 final_adder.U$$212/B
+ sky130_fd_sc_hd__ha_1
XU$$3272 U$$3272/A U$$3287/A VGND VGND VPWR VPWR U$$3272/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$54 _350_/Q _222_/Q VGND VGND VPWR VPWR final_adder.U$$971/B1 final_adder.U$$200/A
+ sky130_fd_sc_hd__ha_1
XU$$3283 U$$3555/B1 U$$3285/A2 U$$3283/B1 U$$3285/B2 VGND VGND VPWR VPWR U$$3284/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$65 _361_/Q _233_/Q VGND VGND VPWR VPWR final_adder.U$$191/B1 final_adder.U$$190/B
+ sky130_fd_sc_hd__ha_1
XFILLER_34_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3294 U$$3294/A1 U$$3320/A2 input65/X U$$3320/B2 VGND VGND VPWR VPWR U$$3295/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$76 _372_/Q _244_/Q VGND VGND VPWR VPWR final_adder.U$$949/B1 final_adder.U$$178/A
+ sky130_fd_sc_hd__ha_1
XU$$2560 U$$3245/A1 U$$2588/A2 U$$3245/B1 U$$2588/B2 VGND VGND VPWR VPWR U$$2561/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$87 _383_/Q _255_/Q VGND VGND VPWR VPWR final_adder.U$$169/B1 final_adder.U$$168/B
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$98 _394_/Q _266_/Q VGND VGND VPWR VPWR final_adder.U$$927/B1 final_adder.U$$156/A
+ sky130_fd_sc_hd__ha_1
XU$$2571 U$$2571/A U$$2577/B VGND VGND VPWR VPWR U$$2571/X sky130_fd_sc_hd__xor2_1
XU$$4409_1781 VGND VGND VPWR VPWR U$$4409_1781/HI U$$4409/B sky130_fd_sc_hd__conb_1
XU$$2582 U$$2582/A1 U$$2588/A2 U$$4502/A1 U$$2588/B2 VGND VGND VPWR VPWR U$$2583/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2593 U$$2593/A U$$2601/B VGND VGND VPWR VPWR U$$2593/X sky130_fd_sc_hd__xor2_1
XFILLER_22_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1870 U$$1870/A U$$1870/B VGND VGND VPWR VPWR U$$1870/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1881 U$$2701/B1 U$$1913/A2 U$$924/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1882/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1892 U$$1892/A U$$1917/A VGND VGND VPWR VPWR U$$1892/X sky130_fd_sc_hd__xor2_1
XFILLER_210_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_89_3 U$$2978/X U$$3111/X U$$3244/X VGND VGND VPWR VPWR dadda_fa_2_90_4/CIN
+ dadda_fa_3_89_0/A sky130_fd_sc_hd__fa_1
XFILLER_192_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_66_2 dadda_fa_4_66_2/A dadda_fa_4_66_2/B dadda_fa_4_66_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_67_0/CIN dadda_fa_5_66_1/CIN sky130_fd_sc_hd__fa_1
XTAP_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_59_1 dadda_fa_4_59_1/A dadda_fa_4_59_1/B dadda_fa_4_59_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/B dadda_fa_5_59_1/B sky130_fd_sc_hd__fa_1
XTAP_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$500 final_adder.U$$500/A final_adder.U$$500/B VGND VGND VPWR VPWR
+ final_adder.U$$616/A sky130_fd_sc_hd__and2_1
XTAP_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$511 final_adder.U$$510/B final_adder.U$$395/X final_adder.U$$387/X
+ VGND VGND VPWR VPWR final_adder.U$$511/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_7_36_0 dadda_fa_7_36_0/A dadda_fa_7_36_0/B dadda_fa_7_36_0/CIN VGND VGND
+ VPWR VPWR _333_/D _204_/D sky130_fd_sc_hd__fa_2
XTAP_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$522 final_adder.U$$530/B final_adder.U$$522/B VGND VGND VPWR VPWR
+ final_adder.U$$642/B sky130_fd_sc_hd__and2_1
XTAP_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$533 final_adder.U$$532/B final_adder.U$$417/X final_adder.U$$409/X
+ VGND VGND VPWR VPWR final_adder.U$$533/X sky130_fd_sc_hd__a21o_1
XTAP_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$544 final_adder.U$$552/B final_adder.U$$544/B VGND VGND VPWR VPWR
+ final_adder.U$$664/B sky130_fd_sc_hd__and2_1
XTAP_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$555 final_adder.U$$554/B final_adder.U$$439/X final_adder.U$$431/X
+ VGND VGND VPWR VPWR final_adder.U$$555/X sky130_fd_sc_hd__a21o_1
XTAP_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$566 final_adder.U$$574/B final_adder.U$$566/B VGND VGND VPWR VPWR
+ final_adder.U$$686/B sky130_fd_sc_hd__and2_1
XTAP_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$405 U$$405/A U$$410/A VGND VGND VPWR VPWR U$$405/X sky130_fd_sc_hd__xor2_1
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater770 U$$366/B2 VGND VGND VPWR VPWR U$$378/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$577 final_adder.U$$576/B final_adder.U$$461/X final_adder.U$$453/X
+ VGND VGND VPWR VPWR final_adder.U$$577/X sky130_fd_sc_hd__a21o_1
XTAP_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$416 U$$414/B U$$410/A U$$412/A U$$411/Y VGND VGND VPWR VPWR U$$416/X sky130_fd_sc_hd__a22o_4
Xrepeater781 U$$2844/B2 VGND VGND VPWR VPWR U$$2828/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$588 final_adder.U$$596/B final_adder.U$$588/B VGND VGND VPWR VPWR
+ final_adder.U$$708/B sky130_fd_sc_hd__and2_1
XU$$427 U$$16/A1 U$$437/A2 U$$703/A1 U$$437/B2 VGND VGND VPWR VPWR U$$428/A sky130_fd_sc_hd__a22o_1
XTAP_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater792 U$$2588/B2 VGND VGND VPWR VPWR U$$2600/B2 sky130_fd_sc_hd__buf_4
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$599 final_adder.U$$598/B final_adder.U$$483/X final_adder.U$$475/X
+ VGND VGND VPWR VPWR final_adder.U$$599/X sky130_fd_sc_hd__a21o_1
XU$$438 U$$438/A U$$474/B VGND VGND VPWR VPWR U$$438/X sky130_fd_sc_hd__xor2_1
XU$$449 U$$38/A1 U$$473/A2 U$$40/A1 U$$473/B2 VGND VGND VPWR VPWR U$$450/A sky130_fd_sc_hd__a22o_1
XFILLER_56_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1305 U$$3389/B VGND VGND VPWR VPWR U$$3395/B sky130_fd_sc_hd__buf_6
Xrepeater1316 U$$3256/B VGND VGND VPWR VPWR U$$3264/B sky130_fd_sc_hd__buf_6
XFILLER_153_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1327 U$$3117/B VGND VGND VPWR VPWR U$$3133/B sky130_fd_sc_hd__buf_8
XFILLER_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1338 input38/X VGND VGND VPWR VPWR U$$3008/B sky130_fd_sc_hd__buf_6
XFILLER_84_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1349 U$$264/B VGND VGND VPWR VPWR U$$218/B sky130_fd_sc_hd__buf_8
XFILLER_101_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_61_1 dadda_fa_3_61_1/A dadda_fa_3_61_1/B dadda_fa_3_61_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_0/CIN dadda_fa_4_61_2/A sky130_fd_sc_hd__fa_1
XFILLER_121_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_54_0 dadda_fa_3_54_0/A dadda_fa_3_54_0/B dadda_fa_3_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_0/B dadda_fa_4_54_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$950 U$$950/A1 U$$950/A2 U$$950/B1 U$$950/B2 VGND VGND VPWR VPWR U$$951/A sky130_fd_sc_hd__a22o_1
XFILLER_211_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1100 U$$1098/Y input8/X U$$962/A U$$1099/X U$$1096/Y VGND VGND VPWR VPWR U$$1100/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_91_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$961 U$$962/A VGND VGND VPWR VPWR U$$961/Y sky130_fd_sc_hd__inv_1
XFILLER_91_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$972 U$$972/A U$$980/B VGND VGND VPWR VPWR U$$972/X sky130_fd_sc_hd__xor2_1
XFILLER_44_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1111 U$$1111/A U$$1139/B VGND VGND VPWR VPWR U$$1111/X sky130_fd_sc_hd__xor2_1
XU$$1122 U$$985/A1 U$$1136/A2 U$$4410/B1 U$$1136/B2 VGND VGND VPWR VPWR U$$1123/A
+ sky130_fd_sc_hd__a22o_1
XU$$983 U$$983/A1 U$$999/A2 U$$983/B1 U$$999/B2 VGND VGND VPWR VPWR U$$984/A sky130_fd_sc_hd__a22o_1
XU$$994 U$$994/A U$$994/B VGND VGND VPWR VPWR U$$994/X sky130_fd_sc_hd__xor2_1
XU$$1133 U$$1133/A U$$1137/B VGND VGND VPWR VPWR U$$1133/X sky130_fd_sc_hd__xor2_1
XFILLER_16_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1144 U$$733/A1 U$$1190/A2 U$$598/A1 U$$1190/B2 VGND VGND VPWR VPWR U$$1145/A sky130_fd_sc_hd__a22o_1
XU$$1155 U$$1155/A U$$1195/B VGND VGND VPWR VPWR U$$1155/X sky130_fd_sc_hd__xor2_1
XFILLER_204_674 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1166 U$$70/A1 U$$1174/A2 U$$2810/B1 U$$1174/B2 VGND VGND VPWR VPWR U$$1167/A sky130_fd_sc_hd__a22o_1
XFILLER_206_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1177 U$$1177/A U$$1223/B VGND VGND VPWR VPWR U$$1177/X sky130_fd_sc_hd__xor2_1
XFILLER_188_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1188 U$$366/A1 U$$1190/A2 U$$94/A1 U$$1190/B2 VGND VGND VPWR VPWR U$$1189/A sky130_fd_sc_hd__a22o_1
XU$$1199 U$$1199/A U$$1205/B VGND VGND VPWR VPWR U$$1199/X sky130_fd_sc_hd__xor2_1
XFILLER_31_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_111_0 dadda_fa_7_111_0/A dadda_fa_7_111_0/B dadda_fa_7_111_0/CIN VGND
+ VGND VPWR VPWR _408_/D _279_/D sky130_fd_sc_hd__fa_1
XFILLER_176_559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_99_2 U$$3264/X U$$3397/X U$$3530/X VGND VGND VPWR VPWR dadda_fa_3_100_1/CIN
+ dadda_fa_3_99_3/B sky130_fd_sc_hd__fa_1
XFILLER_7_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4439_1796 VGND VGND VPWR VPWR U$$4439_1796/HI U$$4439/B sky130_fd_sc_hd__conb_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_76_1 dadda_fa_5_76_1/A dadda_fa_5_76_1/B dadda_fa_5_76_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_77_0/B dadda_fa_7_76_0/A sky130_fd_sc_hd__fa_1
XFILLER_144_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_69_0 dadda_fa_5_69_0/A dadda_fa_5_69_0/B dadda_fa_5_69_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_70_0/A dadda_fa_6_69_0/CIN sky130_fd_sc_hd__fa_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_1_68_8 dadda_fa_1_68_8/A dadda_fa_1_68_8/B dadda_fa_1_68_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_69_3/A dadda_fa_3_68_0/A sky130_fd_sc_hd__fa_1
XFILLER_26_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3080 U$$4450/A1 U$$3082/A2 U$$4452/A1 U$$3082/B2 VGND VGND VPWR VPWR U$$3081/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_8_0 dadda_fa_6_8_0/A dadda_fa_6_8_0/B dadda_fa_6_8_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_9_0/B dadda_fa_7_8_0/CIN sky130_fd_sc_hd__fa_1
XU$$3091 U$$3091/A U$$3117/B VGND VGND VPWR VPWR U$$3091/X sky130_fd_sc_hd__xor2_1
XFILLER_198_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2390 U$$2390/A U$$2426/B VGND VGND VPWR VPWR U$$2390/X sky130_fd_sc_hd__xor2_1
XFILLER_50_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_71_0 dadda_fa_4_71_0/A dadda_fa_4_71_0/B dadda_fa_4_71_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/A dadda_fa_5_71_1/A sky130_fd_sc_hd__fa_1
XFILLER_116_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_87_0 U$$1643/Y U$$1777/X U$$1910/X VGND VGND VPWR VPWR dadda_fa_2_88_3/A
+ dadda_fa_2_87_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_640 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$330 final_adder.U$$332/B final_adder.U$$330/B VGND VGND VPWR VPWR
+ final_adder.U$$456/B sky130_fd_sc_hd__and2_1
XTAP_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$341 final_adder.U$$340/B final_adder.U$$215/X final_adder.U$$213/X
+ VGND VGND VPWR VPWR final_adder.U$$341/X sky130_fd_sc_hd__a21o_1
XTAP_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$352 final_adder.U$$354/B final_adder.U$$352/B VGND VGND VPWR VPWR
+ final_adder.U$$478/B sky130_fd_sc_hd__and2_1
XTAP_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$363 final_adder.U$$362/B final_adder.U$$237/X final_adder.U$$235/X
+ VGND VGND VPWR VPWR final_adder.U$$363/X sky130_fd_sc_hd__a21o_1
XTAP_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$202 U$$202/A U$$212/B VGND VGND VPWR VPWR U$$202/X sky130_fd_sc_hd__xor2_1
XFILLER_206_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$374 final_adder.U$$376/B final_adder.U$$374/B VGND VGND VPWR VPWR
+ final_adder.U$$500/B sky130_fd_sc_hd__and2_1
XTAP_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$213 U$$76/A1 U$$259/A2 U$$78/A1 U$$259/B2 VGND VGND VPWR VPWR U$$214/A sky130_fd_sc_hd__a22o_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$385 final_adder.U$$384/B final_adder.U$$263/X final_adder.U$$259/X
+ VGND VGND VPWR VPWR final_adder.U$$385/X sky130_fd_sc_hd__a21o_1
XTAP_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$224 U$$224/A U$$264/B VGND VGND VPWR VPWR U$$224/X sky130_fd_sc_hd__xor2_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$396 final_adder.U$$400/B final_adder.U$$396/B VGND VGND VPWR VPWR
+ final_adder.U$$520/B sky130_fd_sc_hd__and2_1
XTAP_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$235 U$$98/A1 U$$243/A2 U$$920/B1 U$$243/B2 VGND VGND VPWR VPWR U$$236/A sky130_fd_sc_hd__a22o_1
XU$$246 U$$246/A U$$260/B VGND VGND VPWR VPWR U$$246/X sky130_fd_sc_hd__xor2_1
XTAP_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$257 U$$942/A1 U$$257/A2 U$$944/A1 U$$257/B2 VGND VGND VPWR VPWR U$$258/A sky130_fd_sc_hd__a22o_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$268 U$$268/A U$$272/B VGND VGND VPWR VPWR U$$268/X sky130_fd_sc_hd__xor2_1
XFILLER_60_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$279 U$$277/B U$$274/A U$$275/A U$$274/Y VGND VGND VPWR VPWR U$$279/X sky130_fd_sc_hd__a22o_4
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$7 U$$7/A U$$9/B VGND VGND VPWR VPWR U$$7/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_86_0 dadda_fa_6_86_0/A dadda_fa_6_86_0/B dadda_fa_6_86_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_87_0/B dadda_fa_7_86_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1102 input76/X VGND VGND VPWR VPWR U$$3296/B1 sky130_fd_sc_hd__buf_4
Xrepeater1113 input75/X VGND VGND VPWR VPWR U$$4019/A1 sky130_fd_sc_hd__buf_6
XFILLER_181_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1124 input73/X VGND VGND VPWR VPWR U$$4013/B1 sky130_fd_sc_hd__clkbuf_8
Xrepeater1135 U$$3737/B1 VGND VGND VPWR VPWR U$$860/B1 sky130_fd_sc_hd__buf_4
XFILLER_126_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1146 U$$36/A1 VGND VGND VPWR VPWR U$$719/B1 sky130_fd_sc_hd__buf_6
Xrepeater1157 U$$1084/B VGND VGND VPWR VPWR U$$998/B sky130_fd_sc_hd__buf_6
XFILLER_126_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1168 U$$4144/A1 VGND VGND VPWR VPWR U$$4005/B1 sky130_fd_sc_hd__buf_8
Xrepeater1179 input68/X VGND VGND VPWR VPWR U$$4005/A1 sky130_fd_sc_hd__buf_6
XFILLER_107_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_102_0_1861 VGND VGND VPWR VPWR dadda_fa_2_102_0/A dadda_fa_2_102_0_1861/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_49_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$780 U$$780/A U$$784/B VGND VGND VPWR VPWR U$$780/X sky130_fd_sc_hd__xor2_1
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$791 U$$928/A1 U$$793/A2 U$$930/A1 U$$793/B2 VGND VGND VPWR VPWR U$$792/A sky130_fd_sc_hd__a22o_1
XFILLER_205_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_392 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _255_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_191_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_551 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1680 U$$2425/A1 VGND VGND VPWR VPWR U$$96/A1 sky130_fd_sc_hd__buf_6
Xdadda_fa_1_80_7 U$$3891/X U$$4024/X U$$4157/X VGND VGND VPWR VPWR dadda_fa_2_81_3/A
+ dadda_fa_2_80_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_99_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1691 input102/X VGND VGND VPWR VPWR U$$3245/A1 sky130_fd_sc_hd__buf_6
XFILLER_98_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_73_6 U$$4276/X U$$4409/X input227/X VGND VGND VPWR VPWR dadda_fa_2_74_2/B
+ dadda_fa_2_73_5/B sky130_fd_sc_hd__fa_1
XFILLER_115_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_66_5 input219/X dadda_fa_1_66_5/B dadda_fa_1_66_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_67_2/A dadda_fa_2_66_5/A sky130_fd_sc_hd__fa_2
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_59_4 U$$3184/X U$$3317/X U$$3450/X VGND VGND VPWR VPWR dadda_fa_2_60_1/CIN
+ dadda_fa_2_59_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_29_2 dadda_fa_4_29_2/A dadda_fa_4_29_2/B dadda_fa_4_29_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_30_0/CIN dadda_fa_5_29_1/CIN sky130_fd_sc_hd__fa_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_805 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_979 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1055 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4506 U$$4506/A1 U$$4388/X U$$4508/A1 U$$4512/B2 VGND VGND VPWR VPWR U$$4507/A
+ sky130_fd_sc_hd__a22o_1
XU$$4517 U$$4517/A U$$4517/B VGND VGND VPWR VPWR U$$4517/X sky130_fd_sc_hd__xor2_1
XTAP_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3805 input108/X U$$3819/A2 input110/X U$$3819/B2 VGND VGND VPWR VPWR U$$3806/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_ha_3_18_2 U$$841/X U$$974/X VGND VGND VPWR VPWR dadda_fa_4_19_1/CIN dadda_ha_3_18_2/SUM
+ sky130_fd_sc_hd__ha_1
XTAP_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3816 U$$3816/A U$$3834/B VGND VGND VPWR VPWR U$$3816/X sky130_fd_sc_hd__xor2_1
XTAP_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3827 U$$4099/B1 U$$3833/A2 U$$3829/A1 U$$3833/B2 VGND VGND VPWR VPWR U$$3828/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$160 final_adder.U$$160/A final_adder.U$$160/B VGND VGND VPWR VPWR
+ final_adder.U$$288/B sky130_fd_sc_hd__and2_1
XTAP_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3838 U$$3909/B VGND VGND VPWR VPWR U$$3838/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$171 final_adder.U$$170/B final_adder.U$$941/B1 final_adder.U$$171/B1
+ VGND VGND VPWR VPWR final_adder.U$$171/X sky130_fd_sc_hd__a21o_1
XTAP_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3849 U$$3849/A U$$3879/B VGND VGND VPWR VPWR U$$3849/X sky130_fd_sc_hd__xor2_1
XFILLER_206_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$182 final_adder.U$$182/A final_adder.U$$182/B VGND VGND VPWR VPWR
+ final_adder.U$$310/B sky130_fd_sc_hd__and2_1
XTAP_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_31_2 dadda_fa_3_31_2/A dadda_fa_3_31_2/B dadda_fa_3_31_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_1/A dadda_fa_4_31_2/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$193 final_adder.U$$192/B final_adder.U$$963/B1 final_adder.U$$193/B1
+ VGND VGND VPWR VPWR final_adder.U$$193/X sky130_fd_sc_hd__a21o_1
XTAP_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_24_1 U$$1119/X U$$1252/X U$$1385/X VGND VGND VPWR VPWR dadda_fa_4_25_0/CIN
+ dadda_fa_4_24_2/A sky130_fd_sc_hd__fa_1
XTAP_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_17_0 U$$41/X U$$174/X U$$307/X VGND VGND VPWR VPWR dadda_fa_4_18_1/B dadda_fa_4_17_2/B
+ sky130_fd_sc_hd__fa_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_1143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_387_ _387_/CLK _387_/D VGND VGND VPWR VPWR _387_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_174_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_1114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_83_5 dadda_fa_2_83_5/A dadda_fa_2_83_5/B dadda_fa_2_83_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_84_2/A dadda_fa_4_83_0/A sky130_fd_sc_hd__fa_2
XFILLER_99_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_76_4 dadda_fa_2_76_4/A dadda_fa_2_76_4/B dadda_fa_2_76_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_1/CIN dadda_fa_3_76_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_69_3 dadda_fa_2_69_3/A dadda_fa_2_69_3/B dadda_fa_2_69_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/B dadda_fa_3_69_3/B sky130_fd_sc_hd__fa_1
XFILLER_110_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_922 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_39_1 dadda_fa_5_39_1/A dadda_fa_5_39_1/B dadda_fa_5_39_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_40_0/B dadda_fa_7_39_0/A sky130_fd_sc_hd__fa_2
XFILLER_110_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_977 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_113_1 dadda_fa_5_113_1/A dadda_fa_5_113_1/B dadda_fa_5_113_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_114_0/B dadda_fa_7_113_0/A sky130_fd_sc_hd__fa_1
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_899 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_106_0 dadda_fa_5_106_0/A dadda_fa_5_106_0/B dadda_fa_5_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_107_0/A dadda_fa_6_106_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_191_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_71_3 U$$3341/X U$$3474/X U$$3607/X VGND VGND VPWR VPWR dadda_fa_2_72_1/B
+ dadda_fa_2_71_4/B sky130_fd_sc_hd__fa_1
XFILLER_154_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_64_2 U$$3327/X U$$3460/X U$$3593/X VGND VGND VPWR VPWR dadda_fa_2_65_1/A
+ dadda_fa_2_64_4/A sky130_fd_sc_hd__fa_1
XFILLER_101_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_41_1 dadda_fa_4_41_1/A dadda_fa_4_41_1/B dadda_fa_4_41_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/B dadda_fa_5_41_1/B sky130_fd_sc_hd__fa_1
XFILLER_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_57_1 U$$1584/X U$$1717/X U$$1850/X VGND VGND VPWR VPWR dadda_fa_2_58_0/CIN
+ dadda_fa_2_57_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_34_0 dadda_fa_4_34_0/A dadda_fa_4_34_0/B dadda_fa_4_34_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/A dadda_fa_5_34_1/A sky130_fd_sc_hd__fa_1
XFILLER_28_955 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_476 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ _337_/CLK _310_/D VGND VGND VPWR VPWR _310_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_952 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_241_ _370_/CLK _241_/D VGND VGND VPWR VPWR _241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_172_ _323_/CLK _172_/D VGND VGND VPWR VPWR _172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_86_3 dadda_fa_3_86_3/A dadda_fa_3_86_3/B dadda_fa_3_86_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_87_1/B dadda_fa_4_86_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_79_2 dadda_fa_3_79_2/A dadda_fa_3_79_2/B dadda_fa_3_79_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_1/A dadda_fa_4_79_2/B sky130_fd_sc_hd__fa_1
XFILLER_77_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1017 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_49_0 dadda_fa_6_49_0/A dadda_fa_6_49_0/B dadda_fa_6_49_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_50_0/B dadda_fa_7_49_0/CIN sky130_fd_sc_hd__fa_2
XU$$4303 U$$4440/A1 U$$4381/A2 U$$4440/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4304/A
+ sky130_fd_sc_hd__a22o_1
XU$$4314 U$$4314/A U$$4366/B VGND VGND VPWR VPWR U$$4314/X sky130_fd_sc_hd__xor2_1
XFILLER_133_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4325 input93/X U$$4327/A2 U$$4464/A1 U$$4327/B2 VGND VGND VPWR VPWR U$$4326/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4336 U$$4336/A U$$4354/B VGND VGND VPWR VPWR U$$4336/X sky130_fd_sc_hd__xor2_1
XU$$4347 U$$4484/A1 U$$4361/A2 U$$4484/B1 U$$4361/B2 VGND VGND VPWR VPWR U$$4348/A
+ sky130_fd_sc_hd__a22o_1
XU$$3602 U$$3737/B1 U$$3636/A2 U$$4426/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3603/A
+ sky130_fd_sc_hd__a22o_1
XU$$4358 U$$4358/A input60/X VGND VGND VPWR VPWR U$$4358/X sky130_fd_sc_hd__xor2_1
XU$$3613 U$$3613/A U$$3613/B VGND VGND VPWR VPWR U$$3613/X sky130_fd_sc_hd__xor2_1
XFILLER_203_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3624 U$$3761/A1 U$$3566/X U$$4311/A1 U$$3567/X VGND VGND VPWR VPWR U$$3625/A sky130_fd_sc_hd__a22o_1
XFILLER_18_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4369 U$$4506/A1 U$$4369/A2 U$$4369/B1 U$$4369/B2 VGND VGND VPWR VPWR U$$4370/A
+ sky130_fd_sc_hd__a22o_1
XU$$3635 U$$3635/A U$$3637/B VGND VGND VPWR VPWR U$$3635/X sky130_fd_sc_hd__xor2_1
XU$$2901 U$$709/A1 U$$2919/A2 U$$2901/B1 U$$2919/B2 VGND VGND VPWR VPWR U$$2902/A
+ sky130_fd_sc_hd__a22o_1
XU$$3646 U$$3646/A1 U$$3696/A2 U$$4468/B1 U$$3696/B2 VGND VGND VPWR VPWR U$$3647/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2912 U$$2912/A U$$2920/B VGND VGND VPWR VPWR U$$2912/X sky130_fd_sc_hd__xor2_1
XU$$3657 U$$3657/A U$$3665/B VGND VGND VPWR VPWR U$$3657/X sky130_fd_sc_hd__xor2_1
XU$$3668 input108/X U$$3686/A2 input110/X U$$3686/B2 VGND VGND VPWR VPWR U$$3669/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_108_2 dadda_fa_4_108_2/A dadda_fa_4_108_2/B dadda_fa_4_108_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_109_0/CIN dadda_fa_5_108_1/CIN sky130_fd_sc_hd__fa_1
XU$$2923 U$$3606/B1 U$$2949/A2 U$$3473/A1 U$$2949/B2 VGND VGND VPWR VPWR U$$2924/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3679 U$$3679/A U$$3683/B VGND VGND VPWR VPWR U$$3679/X sky130_fd_sc_hd__xor2_1
XFILLER_19_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2934 U$$2934/A U$$2978/B VGND VGND VPWR VPWR U$$2934/X sky130_fd_sc_hd__xor2_1
XFILLER_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2945 U$$3356/A1 U$$2967/A2 U$$4178/B1 U$$2967/B2 VGND VGND VPWR VPWR U$$2946/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_919 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2956 U$$2956/A U$$3008/B VGND VGND VPWR VPWR U$$2956/X sky130_fd_sc_hd__xor2_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_250 ANTENNA_250/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2967 U$$3102/B1 U$$2967/A2 U$$2967/B1 U$$2967/B2 VGND VGND VPWR VPWR U$$2968/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2978 U$$2978/A U$$2978/B VGND VGND VPWR VPWR U$$2978/X sky130_fd_sc_hd__xor2_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_261 input76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2989 U$$3946/B1 U$$3011/A2 U$$3813/A1 U$$3011/B2 VGND VGND VPWR VPWR U$$2990/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_595 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1083 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_81_2 dadda_fa_2_81_2/A dadda_fa_2_81_2/B dadda_fa_2_81_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/A dadda_fa_3_81_3/A sky130_fd_sc_hd__fa_1
XFILLER_115_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_74_1 dadda_fa_2_74_1/A dadda_fa_2_74_1/B dadda_fa_2_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_0/CIN dadda_fa_3_74_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_114_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_51_0 dadda_fa_5_51_0/A dadda_fa_5_51_0/B dadda_fa_5_51_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_52_0/A dadda_fa_6_51_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_67_0 dadda_fa_2_67_0/A dadda_fa_2_67_0/B dadda_fa_2_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_0/B dadda_fa_3_67_2/B sky130_fd_sc_hd__fa_1
XFILLER_60_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$907 final_adder.U$$136/A final_adder.U$$845/X final_adder.U$$907/B1
+ VGND VGND VPWR VPWR final_adder.U$$907/X sky130_fd_sc_hd__a21o_1
XFILLER_151_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$929 final_adder.U$$158/A final_adder.U$$867/X final_adder.U$$929/B1
+ VGND VGND VPWR VPWR final_adder.U$$929/X sky130_fd_sc_hd__a21o_1
XFILLER_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1040 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_31_clk _255_/CLK VGND VGND VPWR VPWR _414_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_663 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_96_2 dadda_fa_4_96_2/A dadda_fa_4_96_2/B dadda_fa_4_96_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_97_0/CIN dadda_fa_5_96_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_89_1 dadda_fa_4_89_1/A dadda_fa_4_89_1/B dadda_fa_4_89_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/B dadda_fa_5_89_1/B sky130_fd_sc_hd__fa_1
XFILLER_69_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_66_0 dadda_fa_7_66_0/A dadda_fa_7_66_0/B dadda_fa_7_66_0/CIN VGND VGND
+ VPWR VPWR _363_/D _234_/D sky130_fd_sc_hd__fa_1
XFILLER_106_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_1036 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1050 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2208 U$$3987/B1 U$$2226/A2 U$$2621/A1 U$$2226/B2 VGND VGND VPWR VPWR U$$2209/A
+ sky130_fd_sc_hd__a22o_1
XU$$2219 U$$2219/A U$$2273/B VGND VGND VPWR VPWR U$$2219/X sky130_fd_sc_hd__xor2_1
XFILLER_28_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1507 U$$1507/A VGND VGND VPWR VPWR U$$1507/Y sky130_fd_sc_hd__inv_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1518 U$$1518/A U$$1546/B VGND VGND VPWR VPWR U$$1518/X sky130_fd_sc_hd__xor2_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1529 U$$1666/A1 U$$1545/A2 U$$1666/B1 U$$1545/B2 VGND VGND VPWR VPWR U$$1530/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_22_clk _380_/CLK VGND VGND VPWR VPWR _394_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_184_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_224_ _355_/CLK _224_/D VGND VGND VPWR VPWR _224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_91_1 dadda_fa_3_91_1/A dadda_fa_3_91_1/B dadda_fa_3_91_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_0/CIN dadda_fa_4_91_2/A sky130_fd_sc_hd__fa_2
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_84_0 dadda_fa_3_84_0/A dadda_fa_3_84_0/B dadda_fa_3_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_0/B dadda_fa_4_84_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_83_1106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_416 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_394 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater407 U$$624/A2 VGND VGND VPWR VPWR U$$616/A2 sky130_fd_sc_hd__buf_6
Xrepeater418 U$$4369/A2 VGND VGND VPWR VPWR U$$4327/A2 sky130_fd_sc_hd__buf_4
XU$$4100 U$$4100/A U$$4100/B VGND VGND VPWR VPWR U$$4100/X sky130_fd_sc_hd__xor2_1
Xrepeater429 U$$537/A2 VGND VGND VPWR VPWR U$$491/A2 sky130_fd_sc_hd__buf_4
XU$$4111 input57/X VGND VGND VPWR VPWR U$$4113/B sky130_fd_sc_hd__inv_1
XU$$4122 U$$4396/A1 U$$4144/A2 U$$4398/A1 U$$4144/B2 VGND VGND VPWR VPWR U$$4123/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4133 U$$4133/A U$$4165/B VGND VGND VPWR VPWR U$$4133/X sky130_fd_sc_hd__xor2_1
XFILLER_120_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4144 U$$4144/A1 U$$4144/A2 U$$4144/B1 U$$4144/B2 VGND VGND VPWR VPWR U$$4145/A
+ sky130_fd_sc_hd__a22o_1
XU$$3410 U$$3684/A1 U$$3416/A2 U$$3684/B1 U$$3416/B2 VGND VGND VPWR VPWR U$$3411/A
+ sky130_fd_sc_hd__a22o_1
XU$$4155 U$$4155/A U$$4189/B VGND VGND VPWR VPWR U$$4155/X sky130_fd_sc_hd__xor2_1
XU$$3421 U$$3421/A U$$3424/A VGND VGND VPWR VPWR U$$3421/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_113_0 U$$4223/X U$$4356/X U$$4489/X VGND VGND VPWR VPWR dadda_fa_5_114_0/A
+ dadda_fa_5_113_1/A sky130_fd_sc_hd__fa_1
XU$$4166 U$$4440/A1 U$$4176/A2 U$$4440/B1 U$$4176/B2 VGND VGND VPWR VPWR U$$4167/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_46_5 dadda_fa_2_46_5/A dadda_fa_2_46_5/B dadda_fa_2_46_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_47_2/A dadda_fa_4_46_0/A sky130_fd_sc_hd__fa_1
XFILLER_93_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4177 U$$4177/A U$$4243/B VGND VGND VPWR VPWR U$$4177/X sky130_fd_sc_hd__xor2_1
XU$$3432 U$$3432/A U$$3454/B VGND VGND VPWR VPWR U$$3432/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3443 U$$3578/B1 U$$3527/A2 U$$431/A1 U$$3527/B2 VGND VGND VPWR VPWR U$$3444/A
+ sky130_fd_sc_hd__a22o_1
XU$$4188 U$$4323/B1 U$$4188/A2 U$$4188/B1 U$$4188/B2 VGND VGND VPWR VPWR U$$4189/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4199 U$$4199/A U$$4211/B VGND VGND VPWR VPWR U$$4199/X sky130_fd_sc_hd__xor2_1
XFILLER_19_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_39_4 input189/X dadda_fa_2_39_4/B dadda_fa_2_39_4/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_40_1/CIN dadda_fa_3_39_3/CIN sky130_fd_sc_hd__fa_1
XU$$3454 U$$3454/A U$$3454/B VGND VGND VPWR VPWR U$$3454/X sky130_fd_sc_hd__xor2_1
XFILLER_92_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2720 U$$2720/A U$$2739/A VGND VGND VPWR VPWR U$$2720/X sky130_fd_sc_hd__xor2_1
XU$$3465 U$$3737/B1 U$$3503/A2 U$$4426/A1 U$$3503/B2 VGND VGND VPWR VPWR U$$3466/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2731 U$$3414/B1 U$$2735/A2 U$$3281/A1 U$$2735/B2 VGND VGND VPWR VPWR U$$2732/A
+ sky130_fd_sc_hd__a22o_1
XU$$3476 U$$3476/A U$$3480/B VGND VGND VPWR VPWR U$$3476/X sky130_fd_sc_hd__xor2_1
XU$$2742 input36/X VGND VGND VPWR VPWR U$$2742/Y sky130_fd_sc_hd__inv_1
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3487 U$$3761/A1 U$$3489/A2 U$$4311/A1 U$$3489/B2 VGND VGND VPWR VPWR U$$3488/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2753 U$$2753/A U$$2755/B VGND VGND VPWR VPWR U$$2753/X sky130_fd_sc_hd__xor2_1
XU$$3498 U$$3498/A U$$3504/B VGND VGND VPWR VPWR U$$3498/X sky130_fd_sc_hd__xor2_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2764 U$$709/A1 U$$2782/A2 U$$2901/B1 U$$2782/B2 VGND VGND VPWR VPWR U$$2765/A
+ sky130_fd_sc_hd__a22o_1
XU$$2775 U$$2775/A U$$2869/B VGND VGND VPWR VPWR U$$2775/X sky130_fd_sc_hd__xor2_1
XU$$2786 U$$3880/B1 U$$2828/A2 U$$3747/A1 U$$2828/B2 VGND VGND VPWR VPWR U$$2787/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2797 U$$2797/A U$$2797/B VGND VGND VPWR VPWR U$$2797/X sky130_fd_sc_hd__xor2_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_99_0 dadda_fa_5_99_0/A dadda_fa_5_99_0/B dadda_fa_5_99_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_100_0/A dadda_fa_6_99_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_175_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1252 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1088 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$704 final_adder.U$$720/B final_adder.U$$704/B VGND VGND VPWR VPWR
+ final_adder.U$$784/A sky130_fd_sc_hd__and2_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$715 final_adder.U$$714/B final_adder.U$$611/X final_adder.U$$595/X
+ VGND VGND VPWR VPWR final_adder.U$$715/X sky130_fd_sc_hd__a21o_1
XFILLER_69_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_611 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater930 U$$4466/B1 VGND VGND VPWR VPWR U$$4055/B1 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$737 final_adder.U$$720/A final_adder.U$$255/X final_adder.U$$617/X
+ VGND VGND VPWR VPWR final_adder.U$$737/X sky130_fd_sc_hd__a21o_2
Xrepeater941 input95/X VGND VGND VPWR VPWR U$$4466/A1 sky130_fd_sc_hd__buf_6
XFILLER_96_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$748 final_adder.U$$780/B final_adder.U$$748/B VGND VGND VPWR VPWR
+ final_adder.U$$748/X sky130_fd_sc_hd__and2_1
Xrepeater952 U$$4323/B1 VGND VGND VPWR VPWR U$$1448/A1 sky130_fd_sc_hd__buf_6
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$759 final_adder.U$$758/B final_adder.U$$679/X final_adder.U$$647/X
+ VGND VGND VPWR VPWR final_adder.U$$759/X sky130_fd_sc_hd__a21o_1
Xrepeater963 U$$3499/B1 VGND VGND VPWR VPWR U$$896/B1 sky130_fd_sc_hd__buf_4
XFILLER_110_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$609 U$$609/A U$$637/B VGND VGND VPWR VPWR U$$609/X sky130_fd_sc_hd__xor2_1
XFILLER_112_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater974 input91/X VGND VGND VPWR VPWR U$$4458/A1 sky130_fd_sc_hd__buf_6
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_666 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater985 U$$1187/B VGND VGND VPWR VPWR U$$1175/B sky130_fd_sc_hd__buf_6
Xrepeater996 U$$2808/B1 VGND VGND VPWR VPWR U$$892/A1 sky130_fd_sc_hd__buf_4
XFILLER_186_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1509 U$$4375/B1 VGND VGND VPWR VPWR U$$4514/A1 sky130_fd_sc_hd__buf_4
XFILLER_192_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_108_1 U$$3681/X U$$3814/X U$$3947/X VGND VGND VPWR VPWR dadda_fa_4_109_0/CIN
+ dadda_fa_4_108_2/A sky130_fd_sc_hd__fa_1
XFILLER_152_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_362 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4391_1772 VGND VGND VPWR VPWR U$$4391_1772/HI U$$4391/B sky130_fd_sc_hd__conb_1
XFILLER_160_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput290 output290/A VGND VGND VPWR VPWR o[14] sky130_fd_sc_hd__buf_2
XFILLER_43_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4467_1810 VGND VGND VPWR VPWR U$$4467_1810/HI U$$4467/B sky130_fd_sc_hd__conb_1
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_49_3 dadda_fa_3_49_3/A dadda_fa_3_49_3/B dadda_fa_3_49_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_50_1/B dadda_fa_4_49_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2005 U$$2005/A U$$2009/B VGND VGND VPWR VPWR U$$2005/X sky130_fd_sc_hd__xor2_1
XFILLER_74_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2016 U$$2016/A1 U$$2016/A2 U$$2701/B1 U$$2016/B2 VGND VGND VPWR VPWR U$$2017/A
+ sky130_fd_sc_hd__a22o_1
XU$$2027 U$$2027/A U$$2047/B VGND VGND VPWR VPWR U$$2027/X sky130_fd_sc_hd__xor2_1
XU$$2038 U$$940/B1 U$$2040/A2 U$$2312/B1 U$$2040/B2 VGND VGND VPWR VPWR U$$2039/A
+ sky130_fd_sc_hd__a22o_1
XU$$1304 U$$1304/A U$$1316/B VGND VGND VPWR VPWR U$$1304/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2049 U$$2049/A U$$2054/A VGND VGND VPWR VPWR U$$2049/X sky130_fd_sc_hd__xor2_1
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1315 U$$4055/A1 U$$1361/A2 U$$4055/B1 U$$1355/B2 VGND VGND VPWR VPWR U$$1316/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1326 U$$1326/A U$$1330/B VGND VGND VPWR VPWR U$$1326/X sky130_fd_sc_hd__xor2_1
XU$$1337 U$$2842/B1 U$$1337/A2 U$$2709/A1 U$$1337/B2 VGND VGND VPWR VPWR U$$1338/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1348 U$$1348/A input11/X VGND VGND VPWR VPWR U$$1348/X sky130_fd_sc_hd__xor2_1
XFILLER_204_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1359 U$$4236/A1 U$$1361/A2 U$$2318/B1 U$$1367/B2 VGND VGND VPWR VPWR U$$1360/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_399 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_207_ _208_/CLK _207_/D VGND VGND VPWR VPWR _207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1120 final_adder.U$$158/A final_adder.U$$867/X VGND VGND VPWR VPWR
+ output380/A sky130_fd_sc_hd__xor2_1
XFILLER_23_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1131 final_adder.U$$148/B final_adder.U$$919/X VGND VGND VPWR VPWR
+ output265/A sky130_fd_sc_hd__xor2_1
XFILLER_8_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1142 final_adder.U$$136/A final_adder.U$$845/X VGND VGND VPWR VPWR
+ output277/A sky130_fd_sc_hd__xor2_1
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1067 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_2_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _314_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_983 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_51_3 dadda_fa_2_51_3/A dadda_fa_2_51_3/B dadda_fa_2_51_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/B dadda_fa_3_51_3/B sky130_fd_sc_hd__fa_1
XFILLER_61_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_44_2 U$$3075/B input195/X dadda_fa_2_44_2/CIN VGND VGND VPWR VPWR dadda_fa_3_45_1/A
+ dadda_fa_3_44_3/A sky130_fd_sc_hd__fa_1
XFILLER_66_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$11 _307_/Q _179_/Q VGND VGND VPWR VPWR final_adder.U$$245/B1 final_adder.U$$244/B
+ sky130_fd_sc_hd__ha_1
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_21_1 dadda_fa_5_21_1/A dadda_fa_5_21_1/B dadda_fa_5_21_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_22_0/B dadda_fa_7_21_0/A sky130_fd_sc_hd__fa_1
XU$$3240 U$$3240/A U$$3242/B VGND VGND VPWR VPWR U$$3240/X sky130_fd_sc_hd__xor2_1
XFILLER_53_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$22 _318_/Q _190_/Q VGND VGND VPWR VPWR final_adder.U$$233/A2 final_adder.U$$232/A
+ sky130_fd_sc_hd__ha_1
XU$$3251 U$$4484/A1 U$$3255/A2 U$$4484/B1 U$$3255/B2 VGND VGND VPWR VPWR U$$3252/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$33 _329_/Q _201_/Q VGND VGND VPWR VPWR final_adder.U$$223/B1 final_adder.U$$222/B
+ sky130_fd_sc_hd__ha_1
XU$$3262 U$$3262/A U$$3264/B VGND VGND VPWR VPWR U$$3262/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_37_1 U$$1145/X U$$1278/X U$$1411/X VGND VGND VPWR VPWR dadda_fa_3_38_0/CIN
+ dadda_fa_3_37_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_81_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3273 input117/X U$$3277/A2 U$$3684/B1 U$$3277/B2 VGND VGND VPWR VPWR U$$3274/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$44 _340_/Q _212_/Q VGND VGND VPWR VPWR final_adder.U$$981/B1 final_adder.U$$210/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$55 _351_/Q _223_/Q VGND VGND VPWR VPWR final_adder.U$$201/B1 final_adder.U$$200/B
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$66 _362_/Q _234_/Q VGND VGND VPWR VPWR final_adder.U$$959/B1 final_adder.U$$188/A
+ sky130_fd_sc_hd__ha_1
XU$$3284 U$$3284/A U$$3286/B VGND VGND VPWR VPWR U$$3284/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_14_0 dadda_fa_5_14_0/A dadda_fa_5_14_0/B dadda_fa_5_14_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_15_0/A dadda_fa_6_14_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_146_1111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3295 U$$3295/A U$$3321/B VGND VGND VPWR VPWR U$$3295/X sky130_fd_sc_hd__xor2_1
XU$$2550 U$$2550/A1 U$$2600/A2 U$$3922/A1 U$$2600/B2 VGND VGND VPWR VPWR U$$2551/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$77 _373_/Q _245_/Q VGND VGND VPWR VPWR final_adder.U$$179/B1 final_adder.U$$178/B
+ sky130_fd_sc_hd__ha_1
XFILLER_185_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2561 U$$2561/A U$$2603/A VGND VGND VPWR VPWR U$$2561/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$88 _384_/Q _256_/Q VGND VGND VPWR VPWR final_adder.U$$937/B1 final_adder.U$$166/A
+ sky130_fd_sc_hd__ha_1
XU$$2572 U$$2709/A1 U$$2576/A2 U$$2709/B1 U$$2576/B2 VGND VGND VPWR VPWR U$$2573/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$99 _395_/Q _267_/Q VGND VGND VPWR VPWR final_adder.U$$157/B1 final_adder.U$$156/B
+ sky130_fd_sc_hd__ha_1
XFILLER_181_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2583 U$$2583/A U$$2602/A VGND VGND VPWR VPWR U$$2583/X sky130_fd_sc_hd__xor2_1
XU$$2594 U$$3414/B1 U$$2596/A2 U$$3281/A1 U$$2596/B2 VGND VGND VPWR VPWR U$$2595/A
+ sky130_fd_sc_hd__a22o_1
XU$$1860 U$$1860/A U$$1870/B VGND VGND VPWR VPWR U$$1860/X sky130_fd_sc_hd__xor2_1
XFILLER_34_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1871 U$$3102/B1 U$$1877/A2 U$$2967/B1 U$$1877/B2 VGND VGND VPWR VPWR U$$1872/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1882 U$$1882/A U$$1914/B VGND VGND VPWR VPWR U$$1882/X sky130_fd_sc_hd__xor2_1
XU$$1893 U$$2715/A1 U$$1913/A2 U$$2032/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1894/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_40_3 U$$1284/X U$$1417/X VGND VGND VPWR VPWR dadda_fa_2_41_4/CIN dadda_fa_3_40_0/A
+ sky130_fd_sc_hd__ha_1
XTAP_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_59_2 dadda_fa_4_59_2/A dadda_fa_4_59_2/B dadda_fa_4_59_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_60_0/CIN dadda_fa_5_59_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$501 final_adder.U$$500/B final_adder.U$$379/X final_adder.U$$375/X
+ VGND VGND VPWR VPWR final_adder.U$$501/X sky130_fd_sc_hd__a21o_1
XTAP_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$512 final_adder.U$$520/B final_adder.U$$512/B VGND VGND VPWR VPWR
+ final_adder.U$$632/B sky130_fd_sc_hd__and2_1
XTAP_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_313 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$523 final_adder.U$$522/B final_adder.U$$407/X final_adder.U$$399/X
+ VGND VGND VPWR VPWR final_adder.U$$523/X sky130_fd_sc_hd__a21o_1
XTAP_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$534 final_adder.U$$542/B final_adder.U$$534/B VGND VGND VPWR VPWR
+ final_adder.U$$654/B sky130_fd_sc_hd__and2_1
Xdadda_ha_4_10_1 U$$426/X U$$559/X VGND VGND VPWR VPWR dadda_fa_5_11_1/A dadda_ha_4_10_1/SUM
+ sky130_fd_sc_hd__ha_1
XTAP_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$545 final_adder.U$$544/B final_adder.U$$429/X final_adder.U$$421/X
+ VGND VGND VPWR VPWR final_adder.U$$545/X sky130_fd_sc_hd__a21o_1
XTAP_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$556 final_adder.U$$564/B final_adder.U$$556/B VGND VGND VPWR VPWR
+ final_adder.U$$676/B sky130_fd_sc_hd__and2_1
XTAP_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_29_0 dadda_fa_7_29_0/A dadda_fa_7_29_0/B dadda_fa_7_29_0/CIN VGND VGND
+ VPWR VPWR _326_/D _197_/D sky130_fd_sc_hd__fa_2
Xrepeater760 U$$2949/B2 VGND VGND VPWR VPWR U$$2921/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$567 final_adder.U$$566/B final_adder.U$$451/X final_adder.U$$443/X
+ VGND VGND VPWR VPWR final_adder.U$$567/X sky130_fd_sc_hd__a21o_1
XTAP_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$406 U$$678/B1 U$$278/X U$$817/B1 U$$279/X VGND VGND VPWR VPWR U$$407/A sky130_fd_sc_hd__a22o_1
Xrepeater771 U$$394/B2 VGND VGND VPWR VPWR U$$366/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$578 final_adder.U$$586/B final_adder.U$$578/B VGND VGND VPWR VPWR
+ final_adder.U$$698/B sky130_fd_sc_hd__and2_1
XU$$417 U$$417/A1 U$$437/A2 U$$8/A1 U$$437/B2 VGND VGND VPWR VPWR U$$418/A sky130_fd_sc_hd__a22o_1
XTAP_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater782 U$$2745/X VGND VGND VPWR VPWR U$$2844/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$589 final_adder.U$$588/B final_adder.U$$473/X final_adder.U$$465/X
+ VGND VGND VPWR VPWR final_adder.U$$589/X sky130_fd_sc_hd__a21o_1
XU$$428 U$$428/A U$$436/B VGND VGND VPWR VPWR U$$428/X sky130_fd_sc_hd__xor2_1
XFILLER_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater793 U$$2471/X VGND VGND VPWR VPWR U$$2588/B2 sky130_fd_sc_hd__buf_4
XU$$439 U$$850/A1 U$$473/A2 U$$850/B1 U$$473/B2 VGND VGND VPWR VPWR U$$440/A sky130_fd_sc_hd__a22o_1
XFILLER_198_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_703 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4497_1825 VGND VGND VPWR VPWR U$$4497_1825/HI U$$4497/B sky130_fd_sc_hd__conb_1
XFILLER_9_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1252 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1306 U$$3417/B VGND VGND VPWR VPWR U$$3424/A sky130_fd_sc_hd__buf_8
XFILLER_10_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1317 U$$3286/B VGND VGND VPWR VPWR U$$3287/A sky130_fd_sc_hd__buf_6
XFILLER_180_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1328 U$$3117/B VGND VGND VPWR VPWR U$$3083/B sky130_fd_sc_hd__buf_12
XFILLER_158_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1339 U$$2817/B VGND VGND VPWR VPWR U$$2783/B sky130_fd_sc_hd__buf_6
XFILLER_107_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_61_2 dadda_fa_3_61_2/A dadda_fa_3_61_2/B dadda_fa_3_61_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_1/A dadda_fa_4_61_2/B sky130_fd_sc_hd__fa_1
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_780 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_54_1 dadda_fa_3_54_1/A dadda_fa_3_54_1/B dadda_fa_3_54_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_0/CIN dadda_fa_4_54_2/A sky130_fd_sc_hd__fa_1
Xdadda_fa_6_31_0 dadda_fa_6_31_0/A dadda_fa_6_31_0/B dadda_fa_6_31_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_32_0/B dadda_fa_7_31_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_47_0 dadda_fa_3_47_0/A dadda_fa_3_47_0/B dadda_fa_3_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_0/B dadda_fa_4_47_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_169_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$940 U$$940/A1 U$$826/X U$$940/B1 U$$827/X VGND VGND VPWR VPWR U$$941/A sky130_fd_sc_hd__a22o_1
XFILLER_35_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$951 U$$951/A U$$951/B VGND VGND VPWR VPWR U$$951/X sky130_fd_sc_hd__xor2_1
XU$$1101 U$$1099/B input7/X input8/X U$$1096/Y VGND VGND VPWR VPWR U$$1101/X sky130_fd_sc_hd__a22o_4
XU$$962 U$$962/A U$$962/B VGND VGND VPWR VPWR U$$962/X sky130_fd_sc_hd__and2_1
XU$$973 U$$14/A1 U$$979/A2 U$$975/A1 U$$979/B2 VGND VGND VPWR VPWR U$$974/A sky130_fd_sc_hd__a22o_1
XU$$1112 U$$975/A1 U$$1138/A2 U$$18/A1 U$$1138/B2 VGND VGND VPWR VPWR U$$1113/A sky130_fd_sc_hd__a22o_1
XU$$1123 U$$1123/A U$$1137/B VGND VGND VPWR VPWR U$$1123/X sky130_fd_sc_hd__xor2_1
XFILLER_90_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$984 U$$984/A U$$996/B VGND VGND VPWR VPWR U$$984/X sky130_fd_sc_hd__xor2_1
XFILLER_43_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$995 U$$995/A1 U$$999/A2 U$$997/A1 U$$999/B2 VGND VGND VPWR VPWR U$$996/A sky130_fd_sc_hd__a22o_1
XU$$1134 U$$721/B1 U$$1136/A2 U$$999/A1 U$$1136/B2 VGND VGND VPWR VPWR U$$1135/A sky130_fd_sc_hd__a22o_1
XFILLER_71_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1145 U$$1145/A U$$1187/B VGND VGND VPWR VPWR U$$1145/X sky130_fd_sc_hd__xor2_1
XFILLER_91_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_866 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1156 U$$60/A1 U$$1162/A2 U$$62/A1 U$$1162/B2 VGND VGND VPWR VPWR U$$1157/A sky130_fd_sc_hd__a22o_1
XU$$1167 U$$1167/A U$$1175/B VGND VGND VPWR VPWR U$$1167/X sky130_fd_sc_hd__xor2_1
XFILLER_204_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1178 U$$4055/A1 U$$1222/A2 U$$4055/B1 U$$1222/B2 VGND VGND VPWR VPWR U$$1179/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1189 U$$1189/A U$$1209/B VGND VGND VPWR VPWR U$$1189/X sky130_fd_sc_hd__xor2_1
XFILLER_129_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_104_0 dadda_fa_7_104_0/A dadda_fa_7_104_0/B dadda_fa_7_104_0/CIN VGND
+ VGND VPWR VPWR _401_/D _272_/D sky130_fd_sc_hd__fa_1
XFILLER_157_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_99_3 U$$3663/X U$$3796/X U$$3929/X VGND VGND VPWR VPWR dadda_fa_3_100_2/A
+ dadda_fa_3_99_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_5_69_1 dadda_fa_5_69_1/A dadda_fa_5_69_1/B dadda_fa_5_69_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_70_0/B dadda_fa_7_69_0/A sky130_fd_sc_hd__fa_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_411 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3070 U$$3344/A1 U$$3098/A2 U$$3207/B1 U$$3098/B2 VGND VGND VPWR VPWR U$$3071/A
+ sky130_fd_sc_hd__a22o_1
XU$$3081 U$$3081/A U$$3083/B VGND VGND VPWR VPWR U$$3081/X sky130_fd_sc_hd__xor2_1
XU$$3092 U$$4049/B1 U$$3118/A2 U$$3642/A1 U$$3118/B2 VGND VGND VPWR VPWR U$$3093/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2380 U$$2380/A U$$2380/B VGND VGND VPWR VPWR U$$2380/X sky130_fd_sc_hd__xor2_1
XU$$2391 U$$2391/A1 U$$2403/A2 U$$62/B1 U$$2403/B2 VGND VGND VPWR VPWR U$$2392/A sky130_fd_sc_hd__a22o_1
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_555 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1690 U$$594/A1 U$$1736/A2 U$$3473/A1 U$$1736/B2 VGND VGND VPWR VPWR U$$1691/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_71_1 dadda_fa_4_71_1/A dadda_fa_4_71_1/B dadda_fa_4_71_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/B dadda_fa_5_71_1/B sky130_fd_sc_hd__fa_1
XFILLER_104_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_87_1 U$$2043/X U$$2176/X U$$2309/X VGND VGND VPWR VPWR dadda_fa_2_88_3/B
+ dadda_fa_2_87_5/A sky130_fd_sc_hd__fa_1
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_64_0 dadda_fa_4_64_0/A dadda_fa_4_64_0/B dadda_fa_4_64_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/A dadda_fa_5_64_1/A sky130_fd_sc_hd__fa_1
XFILLER_104_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$320 final_adder.U$$322/B final_adder.U$$320/B VGND VGND VPWR VPWR
+ final_adder.U$$446/B sky130_fd_sc_hd__and2_1
XTAP_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$331 final_adder.U$$330/B final_adder.U$$205/X final_adder.U$$203/X
+ VGND VGND VPWR VPWR final_adder.U$$331/X sky130_fd_sc_hd__a21o_1
XTAP_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$342 final_adder.U$$344/B final_adder.U$$342/B VGND VGND VPWR VPWR
+ final_adder.U$$468/B sky130_fd_sc_hd__and2_1
XTAP_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$353 final_adder.U$$352/B final_adder.U$$227/X final_adder.U$$225/X
+ VGND VGND VPWR VPWR final_adder.U$$353/X sky130_fd_sc_hd__a21o_1
XTAP_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$364 final_adder.U$$366/B final_adder.U$$364/B VGND VGND VPWR VPWR
+ final_adder.U$$490/B sky130_fd_sc_hd__and2_1
XTAP_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$203 U$$66/A1 U$$209/A2 U$$68/A1 U$$209/B2 VGND VGND VPWR VPWR U$$204/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$375 final_adder.U$$374/B final_adder.U$$249/X final_adder.U$$247/X
+ VGND VGND VPWR VPWR final_adder.U$$375/X sky130_fd_sc_hd__a21o_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$214 U$$214/A U$$244/B VGND VGND VPWR VPWR U$$214/X sky130_fd_sc_hd__xor2_1
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$386 final_adder.U$$390/B final_adder.U$$386/B VGND VGND VPWR VPWR
+ final_adder.U$$510/B sky130_fd_sc_hd__and2_2
XTAP_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$225 U$$88/A1 U$$263/A2 U$$90/A1 U$$231/B2 VGND VGND VPWR VPWR U$$226/A sky130_fd_sc_hd__a22o_1
XFILLER_55_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater590 U$$1913/A2 VGND VGND VPWR VPWR U$$1915/A2 sky130_fd_sc_hd__buf_8
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$397 final_adder.U$$396/B final_adder.U$$275/X final_adder.U$$271/X
+ VGND VGND VPWR VPWR final_adder.U$$397/X sky130_fd_sc_hd__a21o_1
XFILLER_205_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$236 U$$236/A U$$244/B VGND VGND VPWR VPWR U$$236/X sky130_fd_sc_hd__xor2_1
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$247 U$$521/A1 U$$257/A2 U$$384/B1 U$$257/B2 VGND VGND VPWR VPWR U$$248/A sky130_fd_sc_hd__a22o_1
XTAP_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$258 U$$258/A U$$260/B VGND VGND VPWR VPWR U$$258/X sky130_fd_sc_hd__xor2_1
XU$$269 U$$678/B1 U$$141/X U$$817/B1 U$$142/X VGND VGND VPWR VPWR U$$270/A sky130_fd_sc_hd__a22o_1
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_623 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_526 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$8 U$$8/A1 U$$8/A2 U$$8/B1 U$$8/B2 VGND VGND VPWR VPWR U$$9/A sky130_fd_sc_hd__a22o_1
XFILLER_166_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1103 input76/X VGND VGND VPWR VPWR U$$832/A1 sky130_fd_sc_hd__buf_6
XFILLER_127_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1114 U$$3878/B1 VGND VGND VPWR VPWR U$$864/B1 sky130_fd_sc_hd__buf_4
XFILLER_181_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1125 U$$4289/A1 VGND VGND VPWR VPWR U$$864/A1 sky130_fd_sc_hd__buf_6
Xdadda_ha_0_76_1 U$$1223/X U$$1356/X VGND VGND VPWR VPWR dadda_fa_1_77_8/CIN dadda_fa_2_76_0/A
+ sky130_fd_sc_hd__ha_1
Xrepeater1136 U$$4424/A1 VGND VGND VPWR VPWR U$$3737/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_6_79_0 dadda_fa_6_79_0/A dadda_fa_6_79_0/B dadda_fa_6_79_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_80_0/B dadda_fa_7_79_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater1147 U$$4146/A1 VGND VGND VPWR VPWR U$$36/A1 sky130_fd_sc_hd__buf_4
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1158 U$$1084/B VGND VGND VPWR VPWR U$$968/B sky130_fd_sc_hd__buf_6
XFILLER_181_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_1140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1169 U$$4418/A1 VGND VGND VPWR VPWR U$$4144/A1 sky130_fd_sc_hd__buf_6
XFILLER_4_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_920 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$770 U$$770/A U$$770/B VGND VGND VPWR VPWR U$$770/X sky130_fd_sc_hd__xor2_1
XU$$781 U$$918/A1 U$$783/A2 U$$920/A1 U$$783/B2 VGND VGND VPWR VPWR U$$782/A sky130_fd_sc_hd__a22o_1
XFILLER_91_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$792 U$$792/A U$$794/B VGND VGND VPWR VPWR U$$792/X sky130_fd_sc_hd__xor2_1
XFILLER_90_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_1193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_81_0 dadda_fa_5_81_0/A dadda_fa_5_81_0/B dadda_fa_5_81_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_82_0/A dadda_fa_6_81_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_97_0 U$$2328/Y U$$2462/X U$$2595/X VGND VGND VPWR VPWR dadda_fa_3_98_0/B
+ dadda_fa_3_97_2/B sky130_fd_sc_hd__fa_1
XFILLER_117_468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1670 U$$783/A1 VGND VGND VPWR VPWR U$$920/A1 sky130_fd_sc_hd__buf_4
XFILLER_132_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1681 U$$2425/A1 VGND VGND VPWR VPWR U$$3108/B1 sky130_fd_sc_hd__buf_6
Xrepeater1692 input102/X VGND VGND VPWR VPWR U$$4478/A1 sky130_fd_sc_hd__buf_4
XFILLER_67_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_73_7 dadda_fa_1_73_7/A dadda_fa_1_73_7/B dadda_fa_1_73_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_74_2/CIN dadda_fa_2_73_5/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_66_6 dadda_fa_1_66_6/A dadda_fa_1_66_6/B dadda_fa_1_66_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_2/B dadda_fa_2_66_5/B sky130_fd_sc_hd__fa_1
XFILLER_101_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_59_5 U$$3583/X U$$3716/X U$$3849/X VGND VGND VPWR VPWR dadda_fa_2_60_2/A
+ dadda_fa_2_59_5/A sky130_fd_sc_hd__fa_1
XFILLER_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_7_96_0 dadda_fa_7_96_0/A dadda_fa_7_96_0/B dadda_fa_7_96_0/CIN VGND VGND
+ VPWR VPWR _393_/D _264_/D sky130_fd_sc_hd__fa_1
XFILLER_167_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$4507 U$$4507/A U$$4507/B VGND VGND VPWR VPWR U$$4507/X sky130_fd_sc_hd__xor2_1
XTAP_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_111_0 dadda_fa_6_111_0/A dadda_fa_6_111_0/B dadda_fa_6_111_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_112_0/B dadda_fa_7_111_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3806 U$$3806/A U$$3826/B VGND VGND VPWR VPWR U$$3806/X sky130_fd_sc_hd__xor2_1
XTAP_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3817 U$$3817/A1 U$$3819/A2 input116/X U$$3819/B2 VGND VGND VPWR VPWR U$$3818/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_614 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$150 final_adder.U$$150/A final_adder.U$$150/B VGND VGND VPWR VPWR
+ final_adder.U$$278/B sky130_fd_sc_hd__and2_1
XTAP_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3828 U$$3828/A U$$3834/B VGND VGND VPWR VPWR U$$3828/X sky130_fd_sc_hd__xor2_1
XTAP_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$161 final_adder.U$$160/B final_adder.U$$931/B1 final_adder.U$$161/B1
+ VGND VGND VPWR VPWR final_adder.U$$161/X sky130_fd_sc_hd__a21o_1
XTAP_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$172 final_adder.U$$172/A final_adder.U$$172/B VGND VGND VPWR VPWR
+ final_adder.U$$300/B sky130_fd_sc_hd__and2_1
XTAP_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_422 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3839 U$$3909/B U$$3839/B VGND VGND VPWR VPWR U$$3839/X sky130_fd_sc_hd__and2_1
XTAP_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_31_3 dadda_fa_3_31_3/A dadda_fa_3_31_3/B dadda_fa_3_31_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_32_1/B dadda_fa_4_31_2/CIN sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$183 final_adder.U$$182/B final_adder.U$$953/B1 final_adder.U$$183/B1
+ VGND VGND VPWR VPWR final_adder.U$$183/X sky130_fd_sc_hd__a21o_1
XTAP_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$194 final_adder.U$$194/A final_adder.U$$194/B VGND VGND VPWR VPWR
+ final_adder.U$$322/B sky130_fd_sc_hd__and2_1
XTAP_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_926 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_24_2 U$$1518/X U$$1651/X U$$1679/B VGND VGND VPWR VPWR dadda_fa_4_25_1/A
+ dadda_fa_4_24_2/B sky130_fd_sc_hd__fa_1
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_983 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_386_ _390_/CLK _386_/D VGND VGND VPWR VPWR _386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_76_5 dadda_fa_2_76_5/A dadda_fa_2_76_5/B dadda_fa_2_76_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_77_2/A dadda_fa_4_76_0/A sky130_fd_sc_hd__fa_2
XFILLER_68_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_69_4 dadda_fa_2_69_4/A dadda_fa_2_69_4/B dadda_fa_2_69_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_1/CIN dadda_fa_3_69_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput190 c[3] VGND VGND VPWR VPWR input190/X sky130_fd_sc_hd__buf_4
XFILLER_37_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_106_1 dadda_fa_5_106_1/A dadda_fa_5_106_1/B dadda_fa_5_106_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_107_0/B dadda_fa_7_106_0/A sky130_fd_sc_hd__fa_1
XFILLER_106_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_98_0_1864 VGND VGND VPWR VPWR dadda_fa_2_98_0/A dadda_fa_2_98_0_1864/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_132_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_71_4 U$$3740/X U$$3873/X U$$4006/X VGND VGND VPWR VPWR dadda_fa_2_72_1/CIN
+ dadda_fa_2_71_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_207_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_64_3 U$$3726/X U$$3859/X U$$3992/X VGND VGND VPWR VPWR dadda_fa_2_65_1/B
+ dadda_fa_2_64_4/B sky130_fd_sc_hd__fa_1
XFILLER_101_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_41_2 dadda_fa_4_41_2/A dadda_fa_4_41_2/B dadda_fa_4_41_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_42_0/CIN dadda_fa_5_41_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_57_2 U$$1983/X U$$2116/X U$$2249/X VGND VGND VPWR VPWR dadda_fa_2_58_1/A
+ dadda_fa_2_57_4/A sky130_fd_sc_hd__fa_1
Xdadda_fa_4_34_1 dadda_fa_4_34_1/A dadda_fa_4_34_1/B dadda_fa_4_34_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/B dadda_fa_5_34_1/B sky130_fd_sc_hd__fa_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_11_0 dadda_fa_7_11_0/A dadda_fa_7_11_0/B dadda_fa_7_11_0/CIN VGND VGND
+ VPWR VPWR _308_/D _179_/D sky130_fd_sc_hd__fa_1
XFILLER_43_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_27_0 dadda_fa_4_27_0/A dadda_fa_4_27_0/B dadda_fa_4_27_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/A dadda_fa_5_27_1/A sky130_fd_sc_hd__fa_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_240_ _370_/CLK _240_/D VGND VGND VPWR VPWR _240_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_964 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_171_ _304_/CLK _171_/D VGND VGND VPWR VPWR _171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_0_60_4 U$$1723/X U$$1856/X VGND VGND VPWR VPWR dadda_fa_1_61_7/B dadda_fa_2_60_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_124_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_79_3 dadda_fa_3_79_3/A dadda_fa_3_79_3/B dadda_fa_3_79_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_80_1/B dadda_fa_4_79_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_123_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4304 U$$4304/A U$$4382/B VGND VGND VPWR VPWR U$$4304/X sky130_fd_sc_hd__xor2_1
XU$$4315 U$$4452/A1 U$$4361/A2 input89/X U$$4361/B2 VGND VGND VPWR VPWR U$$4316/A
+ sky130_fd_sc_hd__a22o_1
XU$$4326 U$$4326/A U$$4330/B VGND VGND VPWR VPWR U$$4326/X sky130_fd_sc_hd__xor2_1
XU$$4337 input100/X U$$4349/A2 input101/X U$$4349/B2 VGND VGND VPWR VPWR U$$4338/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_6_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _380_/CLK sky130_fd_sc_hd__clkbuf_8
XU$$4348 U$$4348/A U$$4366/B VGND VGND VPWR VPWR U$$4348/X sky130_fd_sc_hd__xor2_1
XU$$3603 U$$3603/A U$$3637/B VGND VGND VPWR VPWR U$$3603/X sky130_fd_sc_hd__xor2_1
XU$$4359 U$$4496/A1 U$$4361/A2 U$$4498/A1 U$$4361/B2 VGND VGND VPWR VPWR U$$4360/A
+ sky130_fd_sc_hd__a22o_1
XU$$3614 input79/X U$$3644/A2 U$$3614/B1 U$$3644/B2 VGND VGND VPWR VPWR U$$3615/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3625 U$$3625/A input49/X VGND VGND VPWR VPWR U$$3625/X sky130_fd_sc_hd__xor2_1
XU$$3636 U$$3908/B1 U$$3636/A2 U$$3775/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3637/A
+ sky130_fd_sc_hd__a22o_1
XU$$2902 U$$2902/A U$$2920/B VGND VGND VPWR VPWR U$$2902/X sky130_fd_sc_hd__xor2_1
XU$$3647 U$$3647/A U$$3697/B VGND VGND VPWR VPWR U$$3647/X sky130_fd_sc_hd__xor2_1
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2913 U$$4146/A1 U$$2995/A2 input71/X U$$2995/B2 VGND VGND VPWR VPWR U$$2914/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3658 U$$4343/A1 U$$3660/A2 U$$4343/B1 U$$3660/B2 VGND VGND VPWR VPWR U$$3659/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3669 U$$3669/A U$$3698/A VGND VGND VPWR VPWR U$$3669/X sky130_fd_sc_hd__xor2_1
XU$$2924 U$$2924/A U$$2950/B VGND VGND VPWR VPWR U$$2924/X sky130_fd_sc_hd__xor2_1
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_556 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2935 U$$3207/B1 U$$2967/A2 U$$4442/B1 U$$2967/B2 VGND VGND VPWR VPWR U$$2936/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2946 U$$2946/A U$$2968/B VGND VGND VPWR VPWR U$$2946/X sky130_fd_sc_hd__xor2_1
XFILLER_93_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_240 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2957 U$$2957/A1 U$$2967/A2 U$$3368/B1 U$$2967/B2 VGND VGND VPWR VPWR U$$2958/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2968 U$$2968/A U$$2968/B VGND VGND VPWR VPWR U$$2968/X sky130_fd_sc_hd__xor2_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 U$$1/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_262 U$$2967/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2979 U$$3116/A1 U$$2881/X U$$3116/B1 U$$2979/B2 VGND VGND VPWR VPWR U$$2980/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_369_ _370_/CLK _369_/D VGND VGND VPWR VPWR _369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_81_3 dadda_fa_2_81_3/A dadda_fa_2_81_3/B dadda_fa_2_81_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/B dadda_fa_3_81_3/B sky130_fd_sc_hd__fa_1
XFILLER_177_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_74_2 dadda_fa_2_74_2/A dadda_fa_2_74_2/B dadda_fa_2_74_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/A dadda_fa_3_74_3/A sky130_fd_sc_hd__fa_1
XFILLER_25_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_51_1 dadda_fa_5_51_1/A dadda_fa_5_51_1/B dadda_fa_5_51_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_52_0/B dadda_fa_7_51_0/A sky130_fd_sc_hd__fa_1
XFILLER_190_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_67_1 dadda_fa_2_67_1/A dadda_fa_2_67_1/B dadda_fa_2_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_0/CIN dadda_fa_3_67_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_44_0 dadda_fa_5_44_0/A dadda_fa_5_44_0/B dadda_fa_5_44_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_45_0/A dadda_fa_6_44_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_96_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$919 final_adder.U$$148/A final_adder.U$$857/X final_adder.U$$919/B1
+ VGND VGND VPWR VPWR final_adder.U$$919/X sky130_fd_sc_hd__a21o_1
XFILLER_84_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_463 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_723 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_675 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_89_2 dadda_fa_4_89_2/A dadda_fa_4_89_2/B dadda_fa_4_89_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_90_0/CIN dadda_fa_5_89_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_145_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_1048 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_59_0 dadda_fa_7_59_0/A dadda_fa_7_59_0/B dadda_fa_7_59_0/CIN VGND VGND
+ VPWR VPWR _356_/D _227_/D sky130_fd_sc_hd__fa_1
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_62_0 U$$2392/X U$$2525/X U$$2658/X VGND VGND VPWR VPWR dadda_fa_2_63_0/B
+ dadda_fa_2_62_3/B sky130_fd_sc_hd__fa_1
XFILLER_86_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_997 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2209 U$$2209/A U$$2227/B VGND VGND VPWR VPWR U$$2209/X sky130_fd_sc_hd__xor2_1
XFILLER_76_1103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1508 input15/X VGND VGND VPWR VPWR U$$1510/B sky130_fd_sc_hd__inv_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1519 U$$2065/B1 U$$1545/A2 U$$2343/A1 U$$1545/B2 VGND VGND VPWR VPWR U$$1520/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_223_ _355_/CLK _223_/D VGND VGND VPWR VPWR _223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_91_2 dadda_fa_3_91_2/A dadda_fa_3_91_2/B dadda_fa_3_91_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_1/A dadda_fa_4_91_2/B sky130_fd_sc_hd__fa_1
XFILLER_13_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_84_1 dadda_fa_3_84_1/A dadda_fa_3_84_1/B dadda_fa_3_84_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_0/CIN dadda_fa_4_84_2/A sky130_fd_sc_hd__fa_1
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_6_61_0 dadda_fa_6_61_0/A dadda_fa_6_61_0/B dadda_fa_6_61_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_62_0/B dadda_fa_7_61_0/CIN sky130_fd_sc_hd__fa_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_77_0 dadda_fa_3_77_0/A dadda_fa_3_77_0/B dadda_fa_3_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_0/B dadda_fa_4_77_1/CIN sky130_fd_sc_hd__fa_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater408 U$$672/A2 VGND VGND VPWR VPWR U$$624/A2 sky130_fd_sc_hd__buf_4
Xrepeater419 U$$4361/A2 VGND VGND VPWR VPWR U$$4349/A2 sky130_fd_sc_hd__clkbuf_4
XU$$4101 U$$4512/A1 U$$4101/A2 U$$4240/A1 U$$4101/B2 VGND VGND VPWR VPWR U$$4102/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4112 U$$4243/B VGND VGND VPWR VPWR U$$4112/Y sky130_fd_sc_hd__inv_1
XU$$4123 U$$4123/A U$$4145/B VGND VGND VPWR VPWR U$$4123/X sky130_fd_sc_hd__xor2_1
XFILLER_93_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4134 U$$4408/A1 U$$4164/A2 U$$4273/A1 U$$4164/B2 VGND VGND VPWR VPWR U$$4135/A
+ sky130_fd_sc_hd__a22o_1
XU$$3400 U$$3946/B1 U$$3416/A2 U$$251/A1 U$$3416/B2 VGND VGND VPWR VPWR U$$3401/A
+ sky130_fd_sc_hd__a22o_1
XU$$4145 U$$4145/A U$$4145/B VGND VGND VPWR VPWR U$$4145/X sky130_fd_sc_hd__xor2_1
XU$$3411 U$$3411/A U$$3417/B VGND VGND VPWR VPWR U$$3411/X sky130_fd_sc_hd__xor2_1
XU$$4156 input75/X U$$4114/X input77/X U$$4115/X VGND VGND VPWR VPWR U$$4157/A sky130_fd_sc_hd__a22o_1
XU$$3422 input124/X U$$3422/A2 U$$3422/B1 U$$3422/B2 VGND VGND VPWR VPWR U$$3423/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_113_1 input144/X dadda_fa_4_113_1/B dadda_fa_4_113_1/CIN VGND VGND VPWR
+ VPWR dadda_fa_5_114_0/B dadda_fa_5_113_1/B sky130_fd_sc_hd__fa_1
XFILLER_207_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4167 U$$4167/A U$$4246/A VGND VGND VPWR VPWR U$$4167/X sky130_fd_sc_hd__xor2_1
XFILLER_168_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4178 input88/X U$$4188/A2 U$$4178/B1 U$$4188/B2 VGND VGND VPWR VPWR U$$4179/A
+ sky130_fd_sc_hd__a22o_1
XU$$3433 input65/X U$$3453/A2 input76/X U$$3453/B2 VGND VGND VPWR VPWR U$$3434/A sky130_fd_sc_hd__a22o_1
XU$$3444 U$$3444/A U$$3528/B VGND VGND VPWR VPWR U$$3444/X sky130_fd_sc_hd__xor2_1
XU$$4189 U$$4189/A U$$4189/B VGND VGND VPWR VPWR U$$4189/X sky130_fd_sc_hd__xor2_1
XFILLER_81_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2710 U$$2710/A U$$2710/B VGND VGND VPWR VPWR U$$2710/X sky130_fd_sc_hd__xor2_1
XU$$3455 U$$3727/B1 U$$3479/A2 U$$4005/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3456/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_106_0 dadda_fa_4_106_0/A dadda_fa_4_106_0/B dadda_fa_4_106_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/A dadda_fa_5_106_1/A sky130_fd_sc_hd__fa_1
XU$$2721 U$$4228/A1 U$$2737/A2 U$$4365/B1 U$$2737/B2 VGND VGND VPWR VPWR U$$2722/A
+ sky130_fd_sc_hd__a22o_1
XU$$3466 U$$3466/A U$$3504/B VGND VGND VPWR VPWR U$$3466/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_39_5 dadda_fa_2_39_5/A dadda_fa_2_39_5/B dadda_fa_2_39_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_40_2/A dadda_fa_4_39_0/A sky130_fd_sc_hd__fa_1
XFILLER_74_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2732 U$$2732/A U$$2736/B VGND VGND VPWR VPWR U$$2732/X sky130_fd_sc_hd__xor2_1
XFILLER_19_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3477 U$$4162/A1 U$$3479/A2 U$$4027/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3478/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2743 input36/X U$$2743/B VGND VGND VPWR VPWR U$$2743/X sky130_fd_sc_hd__and2_1
XFILLER_73_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3488 U$$3488/A U$$3490/B VGND VGND VPWR VPWR U$$3488/X sky130_fd_sc_hd__xor2_1
XU$$2754 U$$3028/A1 U$$2796/A2 U$$2754/B1 U$$2796/B2 VGND VGND VPWR VPWR U$$2755/A
+ sky130_fd_sc_hd__a22o_1
XU$$3499 U$$3499/A1 U$$3503/A2 U$$3499/B1 U$$3503/B2 VGND VGND VPWR VPWR U$$3500/A
+ sky130_fd_sc_hd__a22o_1
XU$$2765 U$$2765/A U$$2783/B VGND VGND VPWR VPWR U$$2765/X sky130_fd_sc_hd__xor2_1
XU$$2776 U$$4146/A1 U$$2868/A2 input71/X U$$2868/B2 VGND VGND VPWR VPWR U$$2777/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2787 U$$2787/A U$$2817/B VGND VGND VPWR VPWR U$$2787/X sky130_fd_sc_hd__xor2_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2798 U$$4440/B1 U$$2844/A2 U$$4307/A1 U$$2844/B2 VGND VGND VPWR VPWR U$$2799/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_99_1 dadda_fa_5_99_1/A dadda_fa_5_99_1/B dadda_fa_5_99_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_100_0/B dadda_fa_7_99_0/A sky130_fd_sc_hd__fa_1
XFILLER_174_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_864 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1073 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$705 final_adder.U$$704/B final_adder.U$$601/X final_adder.U$$585/X
+ VGND VGND VPWR VPWR final_adder.U$$705/X sky130_fd_sc_hd__a21o_1
XFILLER_68_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$716 final_adder.U$$716/A final_adder.U$$716/B VGND VGND VPWR VPWR
+ final_adder.U$$796/A sky130_fd_sc_hd__and2_1
Xrepeater920 U$$4333/A1 VGND VGND VPWR VPWR U$$3922/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_112_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$727 final_adder.U$$710/A final_adder.U$$623/X final_adder.U$$607/X
+ VGND VGND VPWR VPWR final_adder.U$$727/X sky130_fd_sc_hd__a21o_2
XFILLER_151_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater931 U$$3646/A1 VGND VGND VPWR VPWR U$$3235/A1 sky130_fd_sc_hd__buf_6
XFILLER_69_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater942 input95/X VGND VGND VPWR VPWR U$$3644/A1 sky130_fd_sc_hd__buf_6
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$749 final_adder.U$$748/B final_adder.U$$669/X final_adder.U$$637/X
+ VGND VGND VPWR VPWR final_adder.U$$749/X sky130_fd_sc_hd__a21o_1
Xrepeater953 input93/X VGND VGND VPWR VPWR U$$4323/B1 sky130_fd_sc_hd__buf_4
Xrepeater964 U$$4460/A1 VGND VGND VPWR VPWR U$$3499/B1 sky130_fd_sc_hd__buf_8
Xrepeater975 U$$2949/A1 VGND VGND VPWR VPWR U$$72/A1 sky130_fd_sc_hd__buf_4
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater986 U$$1209/B VGND VGND VPWR VPWR U$$1187/B sky130_fd_sc_hd__buf_8
XFILLER_84_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater997 U$$4178/B1 VGND VGND VPWR VPWR U$$2808/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2189_1728 VGND VGND VPWR VPWR U$$2189_1728/HI U$$2189/B1 sky130_fd_sc_hd__conb_1
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_25 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_4_94_0 dadda_fa_4_94_0/A dadda_fa_4_94_0/B dadda_fa_4_94_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/A dadda_fa_5_94_1/A sky130_fd_sc_hd__fa_1
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_108_2 U$$4080/X U$$4213/X U$$4346/X VGND VGND VPWR VPWR dadda_fa_4_109_1/A
+ dadda_fa_4_108_2/B sky130_fd_sc_hd__fa_1
XFILLER_106_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput280 output280/A VGND VGND VPWR VPWR o[120] sky130_fd_sc_hd__buf_2
XFILLER_121_536 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput291 output291/A VGND VGND VPWR VPWR o[15] sky130_fd_sc_hd__buf_2
XFILLER_43_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2006 U$$2691/A1 U$$2022/A2 U$$2282/A1 U$$2022/B2 VGND VGND VPWR VPWR U$$2007/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_615 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2017 U$$2017/A U$$2017/B VGND VGND VPWR VPWR U$$2017/X sky130_fd_sc_hd__xor2_1
XU$$2028 U$$2165/A1 U$$2052/A2 U$$2715/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2029/A
+ sky130_fd_sc_hd__a22o_1
XU$$2039 U$$2039/A U$$2043/B VGND VGND VPWR VPWR U$$2039/X sky130_fd_sc_hd__xor2_1
XFILLER_204_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1305 U$$72/A1 U$$1311/A2 U$$74/A1 U$$1307/B2 VGND VGND VPWR VPWR U$$1306/A sky130_fd_sc_hd__a22o_1
XU$$1316 U$$1316/A U$$1316/B VGND VGND VPWR VPWR U$$1316/X sky130_fd_sc_hd__xor2_1
XFILLER_128_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1327 U$$94/A1 U$$1337/A2 U$$96/A1 U$$1337/B2 VGND VGND VPWR VPWR U$$1328/A sky130_fd_sc_hd__a22o_1
XU$$1338 U$$1338/A U$$1338/B VGND VGND VPWR VPWR U$$1338/X sky130_fd_sc_hd__xor2_1
XFILLER_31_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1349 U$$527/A1 U$$1353/A2 U$$392/A1 U$$1349/B2 VGND VGND VPWR VPWR U$$1350/A sky130_fd_sc_hd__a22o_1
XFILLER_188_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_206_ _342_/CLK _206_/D VGND VGND VPWR VPWR _206_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1110 final_adder.U$$168/A final_adder.U$$877/X VGND VGND VPWR VPWR
+ output369/A sky130_fd_sc_hd__xor2_1
XFILLER_128_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1121 final_adder.U$$158/B final_adder.U$$929/X VGND VGND VPWR VPWR
+ output381/A sky130_fd_sc_hd__xor2_1
XFILLER_184_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$1132 final_adder.U$$146/A final_adder.U$$855/X VGND VGND VPWR VPWR
+ output266/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1143 final_adder.U$$136/B final_adder.U$$907/X VGND VGND VPWR VPWR
+ output278/A sky130_fd_sc_hd__xor2_1
XFILLER_109_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4515_1834 VGND VGND VPWR VPWR U$$4515_1834/HI U$$4515/B sky130_fd_sc_hd__conb_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1079 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_51_4 dadda_fa_2_51_4/A dadda_fa_2_51_4/B dadda_fa_2_51_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_1/CIN dadda_fa_3_51_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_44_3 dadda_fa_2_44_3/A dadda_fa_2_44_3/B dadda_fa_2_44_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_1/B dadda_fa_3_44_3/B sky130_fd_sc_hd__fa_2
XFILLER_54_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3230 U$$3230/A U$$3244/B VGND VGND VPWR VPWR U$$3230/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$12 _308_/Q _180_/Q VGND VGND VPWR VPWR final_adder.U$$243/A2 final_adder.U$$242/A
+ sky130_fd_sc_hd__ha_1
XU$$3241 U$$3378/A1 U$$3241/A2 U$$3243/A1 U$$3241/B2 VGND VGND VPWR VPWR U$$3242/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$23 _319_/Q _191_/Q VGND VGND VPWR VPWR final_adder.U$$233/B1 final_adder.U$$232/B
+ sky130_fd_sc_hd__ha_1
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$34 _330_/Q _202_/Q VGND VGND VPWR VPWR final_adder.U$$991/B1 final_adder.U$$220/A
+ sky130_fd_sc_hd__ha_1
XU$$3252 U$$3252/A U$$3256/B VGND VGND VPWR VPWR U$$3252/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_37_2 U$$1544/X U$$1677/X U$$1810/X VGND VGND VPWR VPWR dadda_fa_3_38_1/A
+ dadda_fa_3_37_3/A sky130_fd_sc_hd__fa_1
XU$$3263 U$$384/B1 U$$3263/A2 U$$251/A1 U$$3263/B2 VGND VGND VPWR VPWR U$$3264/A sky130_fd_sc_hd__a22o_1
XU$$3274 U$$3274/A U$$3287/A VGND VGND VPWR VPWR U$$3274/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$45 _341_/Q _213_/Q VGND VGND VPWR VPWR final_adder.U$$211/B1 final_adder.U$$210/B
+ sky130_fd_sc_hd__ha_1
XFILLER_59_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$56 _352_/Q _224_/Q VGND VGND VPWR VPWR final_adder.U$$969/B1 final_adder.U$$198/A
+ sky130_fd_sc_hd__ha_1
XU$$3285 U$$3557/B1 U$$3285/A2 U$$3285/B1 U$$3285/B2 VGND VGND VPWR VPWR U$$3286/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2540 U$$3499/A1 U$$2470/X U$$3499/B1 U$$2471/X VGND VGND VPWR VPWR U$$2541/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$67 _363_/Q _235_/Q VGND VGND VPWR VPWR final_adder.U$$189/B1 final_adder.U$$188/B
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_5_14_1 dadda_fa_5_14_1/A dadda_fa_5_14_1/B dadda_fa_5_14_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_15_0/B dadda_fa_7_14_0/A sky130_fd_sc_hd__fa_1
XU$$2551 U$$2551/A U$$2601/B VGND VGND VPWR VPWR U$$2551/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$78 _374_/Q _246_/Q VGND VGND VPWR VPWR final_adder.U$$947/B1 final_adder.U$$176/A
+ sky130_fd_sc_hd__ha_1
XFILLER_185_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3296 input65/X U$$3320/A2 U$$3296/B1 U$$3320/B2 VGND VGND VPWR VPWR U$$3297/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2562 U$$3245/B1 U$$2470/X U$$3112/A1 U$$2471/X VGND VGND VPWR VPWR U$$2563/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$89 _385_/Q _257_/Q VGND VGND VPWR VPWR final_adder.U$$167/B1 final_adder.U$$166/B
+ sky130_fd_sc_hd__ha_1
XFILLER_179_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2573 U$$2573/A U$$2577/B VGND VGND VPWR VPWR U$$2573/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2584 U$$4228/A1 U$$2588/A2 U$$4365/B1 U$$2588/B2 VGND VGND VPWR VPWR U$$2585/A
+ sky130_fd_sc_hd__a22o_1
XU$$2595 U$$2595/A U$$2597/B VGND VGND VPWR VPWR U$$2595/X sky130_fd_sc_hd__xor2_1
XFILLER_146_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1850 U$$1850/A U$$1917/A VGND VGND VPWR VPWR U$$1850/X sky130_fd_sc_hd__xor2_1
XU$$1861 U$$763/B1 U$$1869/A2 U$$630/A1 U$$1869/B2 VGND VGND VPWR VPWR U$$1862/A sky130_fd_sc_hd__a22o_1
XU$$1872 U$$1872/A U$$1878/B VGND VGND VPWR VPWR U$$1872/X sky130_fd_sc_hd__xor2_1
XFILLER_21_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1883 U$$924/A1 U$$1913/A2 U$$789/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1884/A sky130_fd_sc_hd__a22o_1
XFILLER_210_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1894 U$$1894/A U$$1914/B VGND VGND VPWR VPWR U$$1894/X sky130_fd_sc_hd__xor2_1
XFILLER_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_159_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_831 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1084 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_623 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$513 final_adder.U$$512/B final_adder.U$$397/X final_adder.U$$389/X
+ VGND VGND VPWR VPWR final_adder.U$$513/X sky130_fd_sc_hd__a21o_1
XTAP_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$524 final_adder.U$$532/B final_adder.U$$524/B VGND VGND VPWR VPWR
+ final_adder.U$$644/B sky130_fd_sc_hd__and2_1
XFILLER_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$535 final_adder.U$$534/B final_adder.U$$419/X final_adder.U$$411/X
+ VGND VGND VPWR VPWR final_adder.U$$535/X sky130_fd_sc_hd__a21o_1
XTAP_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$546 final_adder.U$$554/B final_adder.U$$546/B VGND VGND VPWR VPWR
+ final_adder.U$$666/B sky130_fd_sc_hd__and2_1
XTAP_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater750 U$$3098/B2 VGND VGND VPWR VPWR U$$3060/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$557 final_adder.U$$556/B final_adder.U$$441/X final_adder.U$$433/X
+ VGND VGND VPWR VPWR final_adder.U$$557/X sky130_fd_sc_hd__a21o_1
XTAP_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater761 U$$2949/B2 VGND VGND VPWR VPWR U$$2919/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$568 final_adder.U$$576/B final_adder.U$$568/B VGND VGND VPWR VPWR
+ final_adder.U$$688/B sky130_fd_sc_hd__and2_1
XTAP_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater772 U$$279/X VGND VGND VPWR VPWR U$$394/B2 sky130_fd_sc_hd__buf_6
XU$$407 U$$407/A U$$410/A VGND VGND VPWR VPWR U$$407/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$579 final_adder.U$$578/B final_adder.U$$463/X final_adder.U$$455/X
+ VGND VGND VPWR VPWR final_adder.U$$579/X sky130_fd_sc_hd__a21o_1
XU$$418 U$$418/A U$$436/B VGND VGND VPWR VPWR U$$418/X sky130_fd_sc_hd__xor2_1
Xrepeater783 U$$2683/B2 VGND VGND VPWR VPWR U$$2625/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_85_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$429 U$$703/A1 U$$515/A2 U$$431/A1 U$$515/B2 VGND VGND VPWR VPWR U$$430/A sky130_fd_sc_hd__a22o_1
XFILLER_38_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater794 U$$2524/B2 VGND VGND VPWR VPWR U$$2490/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_204_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1307 U$$3389/B VGND VGND VPWR VPWR U$$3417/B sky130_fd_sc_hd__buf_8
XFILLER_197_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_113_0 U$$3424/Y U$$3558/X U$$3691/X VGND VGND VPWR VPWR dadda_fa_4_114_1/CIN
+ dadda_fa_4_113_2/B sky130_fd_sc_hd__fa_1
XFILLER_165_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1318 U$$3256/B VGND VGND VPWR VPWR U$$3286/B sky130_fd_sc_hd__buf_6
XFILLER_181_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1329 U$$3151/A VGND VGND VPWR VPWR U$$3117/B sky130_fd_sc_hd__buf_6
XFILLER_107_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_83 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_61_3 dadda_fa_3_61_3/A dadda_fa_3_61_3/B dadda_fa_3_61_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_62_1/B dadda_fa_4_61_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_95_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$271_1736 VGND VGND VPWR VPWR U$$271_1736/HI U$$271/B1 sky130_fd_sc_hd__conb_1
XFILLER_94_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_54_2 dadda_fa_3_54_2/A dadda_fa_3_54_2/B dadda_fa_3_54_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_1/A dadda_fa_4_54_2/B sky130_fd_sc_hd__fa_1
XFILLER_85_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_47_1 dadda_fa_3_47_1/A dadda_fa_3_47_1/B dadda_fa_3_47_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_0/CIN dadda_fa_4_47_2/A sky130_fd_sc_hd__fa_1
XFILLER_63_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_24_0 dadda_fa_6_24_0/A dadda_fa_6_24_0/B dadda_fa_6_24_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_25_0/B dadda_fa_7_24_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$930 U$$930/A1 U$$938/A2 U$$930/B1 U$$938/B2 VGND VGND VPWR VPWR U$$931/A sky130_fd_sc_hd__a22o_1
XU$$941 U$$941/A U$$959/A VGND VGND VPWR VPWR U$$941/X sky130_fd_sc_hd__xor2_1
XFILLER_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$952 U$$952/A1 U$$826/X U$$954/A1 U$$827/X VGND VGND VPWR VPWR U$$953/A sky130_fd_sc_hd__a22o_1
XU$$1102 U$$1102/A1 U$$1138/A2 U$$967/A1 U$$1138/B2 VGND VGND VPWR VPWR U$$1103/A
+ sky130_fd_sc_hd__a22o_1
XU$$963 U$$961/Y input6/X input5/X U$$962/X U$$959/Y VGND VGND VPWR VPWR U$$963/X
+ sky130_fd_sc_hd__a32o_4
XU$$974 U$$974/A U$$980/B VGND VGND VPWR VPWR U$$974/X sky130_fd_sc_hd__xor2_1
XU$$1113 U$$1113/A U$$1139/B VGND VGND VPWR VPWR U$$1113/X sky130_fd_sc_hd__xor2_1
XFILLER_62_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1124 U$$2220/A1 U$$1162/A2 U$$989/A1 U$$1162/B2 VGND VGND VPWR VPWR U$$1125/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$985 U$$985/A1 U$$999/A2 U$$987/A1 U$$999/B2 VGND VGND VPWR VPWR U$$986/A sky130_fd_sc_hd__a22o_1
XFILLER_204_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$996 U$$996/A U$$996/B VGND VGND VPWR VPWR U$$996/X sky130_fd_sc_hd__xor2_1
XFILLER_90_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1135 U$$1135/A U$$1137/B VGND VGND VPWR VPWR U$$1135/X sky130_fd_sc_hd__xor2_1
XU$$1146 U$$598/A1 U$$1190/A2 U$$598/B1 U$$1190/B2 VGND VGND VPWR VPWR U$$1147/A sky130_fd_sc_hd__a22o_1
XFILLER_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1157 U$$1157/A U$$1195/B VGND VGND VPWR VPWR U$$1157/X sky130_fd_sc_hd__xor2_1
XFILLER_71_692 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_3_112_2 U$$4088/X U$$4221/X VGND VGND VPWR VPWR dadda_fa_4_113_2/A dadda_ha_3_112_2/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_149_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1168 U$$72/A1 U$$1174/A2 U$$74/A1 U$$1174/B2 VGND VGND VPWR VPWR U$$1169/A sky130_fd_sc_hd__a22o_1
XU$$1179 U$$1179/A U$$1223/B VGND VGND VPWR VPWR U$$1179/X sky130_fd_sc_hd__xor2_1
XFILLER_204_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1097 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_99_4 U$$4062/X U$$4195/X U$$4328/X VGND VGND VPWR VPWR dadda_fa_3_100_2/B
+ dadda_fa_4_99_0/A sky130_fd_sc_hd__fa_1
XFILLER_171_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_447 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_42_0 U$$1953/X U$$2086/X U$$2219/X VGND VGND VPWR VPWR dadda_fa_3_43_0/B
+ dadda_fa_3_42_2/B sky130_fd_sc_hd__fa_1
XFILLER_39_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3060 U$$3606/B1 U$$3060/A2 U$$3473/A1 U$$3060/B2 VGND VGND VPWR VPWR U$$3061/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3071 U$$3071/A U$$3077/B VGND VGND VPWR VPWR U$$3071/X sky130_fd_sc_hd__xor2_1
XU$$3082 U$$4452/A1 U$$3082/A2 U$$4454/A1 U$$3082/B2 VGND VGND VPWR VPWR U$$3083/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3093 U$$3093/A U$$3117/B VGND VGND VPWR VPWR U$$3093/X sky130_fd_sc_hd__xor2_1
XU$$2370 U$$2370/A U$$2380/B VGND VGND VPWR VPWR U$$2370/X sky130_fd_sc_hd__xor2_1
XFILLER_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2381 U$$3749/B1 U$$2459/A2 input80/X U$$2459/B2 VGND VGND VPWR VPWR U$$2382/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2392 U$$2392/A U$$2442/B VGND VGND VPWR VPWR U$$2392/X sky130_fd_sc_hd__xor2_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1680 U$$993/B1 U$$1688/A2 U$$997/A1 U$$1688/B2 VGND VGND VPWR VPWR U$$1681/A sky130_fd_sc_hd__a22o_1
XFILLER_179_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_528 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1691 U$$1691/A U$$1739/B VGND VGND VPWR VPWR U$$1691/X sky130_fd_sc_hd__xor2_1
XFILLER_33_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_1_88_4 U$$3242/X U$$3375/X VGND VGND VPWR VPWR dadda_fa_2_89_4/CIN dadda_fa_3_88_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_71_2 dadda_fa_4_71_2/A dadda_fa_4_71_2/B dadda_fa_4_71_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_72_0/CIN dadda_fa_5_71_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_87_2 U$$2442/X U$$2575/X U$$2708/X VGND VGND VPWR VPWR dadda_fa_2_88_3/CIN
+ dadda_fa_2_87_5/B sky130_fd_sc_hd__fa_1
XFILLER_104_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_64_1 dadda_fa_4_64_1/A dadda_fa_4_64_1/B dadda_fa_4_64_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/B dadda_fa_5_64_1/B sky130_fd_sc_hd__fa_1
XFILLER_118_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_41_0 dadda_fa_7_41_0/A dadda_fa_7_41_0/B dadda_fa_7_41_0/CIN VGND VGND
+ VPWR VPWR _338_/D _209_/D sky130_fd_sc_hd__fa_2
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_57_0 dadda_fa_4_57_0/A dadda_fa_4_57_0/B dadda_fa_4_57_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/A dadda_fa_5_57_1/A sky130_fd_sc_hd__fa_1
XTAP_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$310 final_adder.U$$312/B final_adder.U$$310/B VGND VGND VPWR VPWR
+ final_adder.U$$436/B sky130_fd_sc_hd__and2_1
XTAP_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$321 final_adder.U$$320/B final_adder.U$$195/X final_adder.U$$193/X
+ VGND VGND VPWR VPWR final_adder.U$$321/X sky130_fd_sc_hd__a21o_1
XFILLER_131_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$332 final_adder.U$$334/B final_adder.U$$332/B VGND VGND VPWR VPWR
+ final_adder.U$$458/B sky130_fd_sc_hd__and2_1
XTAP_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$343 final_adder.U$$342/B final_adder.U$$217/X final_adder.U$$215/X
+ VGND VGND VPWR VPWR final_adder.U$$343/X sky130_fd_sc_hd__a21o_1
XTAP_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$354 final_adder.U$$356/B final_adder.U$$354/B VGND VGND VPWR VPWR
+ final_adder.U$$480/B sky130_fd_sc_hd__and2_1
XTAP_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$365 final_adder.U$$364/B final_adder.U$$239/X final_adder.U$$237/X
+ VGND VGND VPWR VPWR final_adder.U$$365/X sky130_fd_sc_hd__a21o_1
XTAP_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$204 U$$204/A U$$212/B VGND VGND VPWR VPWR U$$204/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$376 final_adder.U$$378/B final_adder.U$$376/B VGND VGND VPWR VPWR
+ final_adder.U$$498/A sky130_fd_sc_hd__and2_1
XTAP_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$215 U$$78/A1 U$$217/A2 U$$80/A1 U$$217/B2 VGND VGND VPWR VPWR U$$216/A sky130_fd_sc_hd__a22o_1
Xrepeater580 U$$2046/A2 VGND VGND VPWR VPWR U$$2052/A2 sky130_fd_sc_hd__buf_6
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$387 final_adder.U$$386/B final_adder.U$$265/X final_adder.U$$261/X
+ VGND VGND VPWR VPWR final_adder.U$$387/X sky130_fd_sc_hd__a21o_1
XTAP_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$226 U$$226/A U$$264/B VGND VGND VPWR VPWR U$$226/X sky130_fd_sc_hd__xor2_1
Xrepeater591 U$$1785/X VGND VGND VPWR VPWR U$$1913/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$398 final_adder.U$$402/B final_adder.U$$398/B VGND VGND VPWR VPWR
+ final_adder.U$$522/B sky130_fd_sc_hd__and2_1
XTAP_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$237 U$$920/B1 U$$243/A2 U$$787/A1 U$$243/B2 VGND VGND VPWR VPWR U$$238/A sky130_fd_sc_hd__a22o_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$248 U$$248/A U$$260/B VGND VGND VPWR VPWR U$$248/X sky130_fd_sc_hd__xor2_1
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$259 U$$944/A1 U$$259/A2 U$$944/B1 U$$259/B2 VGND VGND VPWR VPWR U$$260/A sky130_fd_sc_hd__a22o_1
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$9 U$$9/A U$$9/B VGND VGND VPWR VPWR U$$9/X sky130_fd_sc_hd__xor2_1
XFILLER_166_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1104 U$$4394/A1 VGND VGND VPWR VPWR U$$3159/B1 sky130_fd_sc_hd__buf_6
Xrepeater1115 U$$3058/A1 VGND VGND VPWR VPWR U$$727/B1 sky130_fd_sc_hd__buf_4
Xrepeater1126 U$$3876/B1 VGND VGND VPWR VPWR U$$727/A1 sky130_fd_sc_hd__buf_4
Xrepeater1137 input72/X VGND VGND VPWR VPWR U$$4424/A1 sky130_fd_sc_hd__buf_6
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1148 U$$995/A1 VGND VGND VPWR VPWR U$$993/B1 sky130_fd_sc_hd__buf_6
Xrepeater1159 U$$1076/B VGND VGND VPWR VPWR U$$1084/B sky130_fd_sc_hd__buf_12
XFILLER_113_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_75_0 U$$821/Y U$$955/X U$$1088/X VGND VGND VPWR VPWR dadda_fa_1_76_8/A
+ dadda_fa_1_75_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_171_1068 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$760 U$$760/A U$$796/B VGND VGND VPWR VPWR U$$760/X sky130_fd_sc_hd__xor2_1
XFILLER_90_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$771 U$$84/B1 U$$783/A2 U$$910/A1 U$$783/B2 VGND VGND VPWR VPWR U$$772/A sky130_fd_sc_hd__a22o_1
XU$$782 U$$782/A U$$784/B VGND VGND VPWR VPWR U$$782/X sky130_fd_sc_hd__xor2_1
XFILLER_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$793 U$$930/A1 U$$793/A2 U$$930/B1 U$$793/B2 VGND VGND VPWR VPWR U$$794/A sky130_fd_sc_hd__a22o_1
XFILLER_188_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_5_81_1 dadda_fa_5_81_1/A dadda_fa_5_81_1/B dadda_fa_5_81_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_82_0/B dadda_fa_7_81_0/A sky130_fd_sc_hd__fa_2
XFILLER_144_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_97_1 U$$2728/X U$$2861/X U$$2994/X VGND VGND VPWR VPWR dadda_fa_3_98_0/CIN
+ dadda_fa_3_97_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_145_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_74_0 dadda_fa_5_74_0/A dadda_fa_5_74_0/B dadda_fa_5_74_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_75_0/A dadda_fa_6_74_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_126_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1660 input106/X VGND VGND VPWR VPWR U$$4484/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_99_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1671 U$$2016/A1 VGND VGND VPWR VPWR U$$98/A1 sky130_fd_sc_hd__buf_6
XFILLER_193_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1682 U$$3245/B1 VGND VGND VPWR VPWR U$$2425/A1 sky130_fd_sc_hd__buf_6
XFILLER_116_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1693 input101/X VGND VGND VPWR VPWR U$$4476/A1 sky130_fd_sc_hd__buf_4
XFILLER_63_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_73_8 dadda_fa_1_73_8/A dadda_fa_1_73_8/B dadda_fa_1_73_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_74_3/A dadda_fa_3_73_0/A sky130_fd_sc_hd__fa_1
XFILLER_99_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_66_7 dadda_fa_1_66_7/A dadda_fa_1_66_7/B dadda_fa_1_66_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_2/CIN dadda_fa_2_66_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_6_1054 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_59_6 U$$3982/X input211/X dadda_fa_1_59_6/CIN VGND VGND VPWR VPWR dadda_fa_2_60_2/B
+ dadda_fa_2_59_5/B sky130_fd_sc_hd__fa_1
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_924 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_89_0 dadda_fa_7_89_0/A dadda_fa_7_89_0/B dadda_fa_7_89_0/CIN VGND VGND
+ VPWR VPWR _386_/D _257_/D sky130_fd_sc_hd__fa_2
XFILLER_163_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_1155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_92_0 dadda_fa_1_92_0/A U$$2053/X U$$2186/X VGND VGND VPWR VPWR dadda_fa_2_93_4/CIN
+ dadda_fa_2_92_5/B sky130_fd_sc_hd__fa_1
XFILLER_190_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4508 U$$4508/A1 U$$4388/X U$$4510/A1 U$$4512/B2 VGND VGND VPWR VPWR U$$4509/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$140 final_adder.U$$140/A final_adder.U$$140/B VGND VGND VPWR VPWR
+ final_adder.U$$268/B sky130_fd_sc_hd__and2_1
XU$$3807 U$$3944/A1 U$$3819/A2 U$$3944/B1 U$$3819/B2 VGND VGND VPWR VPWR U$$3808/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3818 U$$3818/A U$$3826/B VGND VGND VPWR VPWR U$$3818/X sky130_fd_sc_hd__xor2_1
XFILLER_57_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$151 final_adder.U$$150/B final_adder.U$$921/B1 final_adder.U$$151/B1
+ VGND VGND VPWR VPWR final_adder.U$$151/X sky130_fd_sc_hd__a21o_1
XTAP_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3829 U$$3829/A1 U$$3833/A2 U$$4103/B1 U$$3833/B2 VGND VGND VPWR VPWR U$$3830/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$162 final_adder.U$$162/A final_adder.U$$162/B VGND VGND VPWR VPWR
+ final_adder.U$$290/B sky130_fd_sc_hd__and2_1
Xdadda_fa_6_104_0 dadda_fa_6_104_0/A dadda_fa_6_104_0/B dadda_fa_6_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_105_0/B dadda_fa_7_104_0/CIN sky130_fd_sc_hd__fa_2
XTAP_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$173 final_adder.U$$172/B final_adder.U$$943/B1 final_adder.U$$173/B1
+ VGND VGND VPWR VPWR final_adder.U$$173/X sky130_fd_sc_hd__a21o_1
XTAP_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$184 final_adder.U$$184/A final_adder.U$$184/B VGND VGND VPWR VPWR
+ final_adder.U$$312/B sky130_fd_sc_hd__and2_1
XTAP_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_968 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$195 final_adder.U$$194/B final_adder.U$$965/B1 final_adder.U$$195/B1
+ VGND VGND VPWR VPWR final_adder.U$$195/X sky130_fd_sc_hd__a21o_1
XFILLER_166_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_24_3 input173/X dadda_fa_3_24_3/B dadda_fa_3_24_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_25_1/B dadda_fa_4_24_2/CIN sky130_fd_sc_hd__fa_1
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_995 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_385_ _385_/CLK _385_/D VGND VGND VPWR VPWR _385_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_91_0 dadda_fa_6_91_0/A dadda_fa_6_91_0/B dadda_fa_6_91_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_92_0/B dadda_fa_7_91_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_103_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_69_5 dadda_fa_2_69_5/A dadda_fa_2_69_5/B dadda_fa_2_69_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_70_2/A dadda_fa_4_69_0/A sky130_fd_sc_hd__fa_1
XFILLER_23_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput180 c[30] VGND VGND VPWR VPWR input180/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput191 c[40] VGND VGND VPWR VPWR input191/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_1158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$590 U$$727/A1 U$$624/A2 U$$727/B1 U$$624/B2 VGND VGND VPWR VPWR U$$591/A sky130_fd_sc_hd__a22o_1
XFILLER_211_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_884 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1490 U$$956/A1 VGND VGND VPWR VPWR U$$1504/A1 sky130_fd_sc_hd__buf_6
XFILLER_28_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1044 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_71_5 U$$4139/X U$$4272/X U$$4405/X VGND VGND VPWR VPWR dadda_fa_2_72_2/A
+ dadda_fa_2_71_5/A sky130_fd_sc_hd__fa_1
XFILLER_8_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_857 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_4 U$$4125/X U$$4258/X U$$4391/X VGND VGND VPWR VPWR dadda_fa_2_65_1/CIN
+ dadda_fa_2_64_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_57_3 U$$2382/X U$$2515/X U$$2648/X VGND VGND VPWR VPWR dadda_fa_2_58_1/B
+ dadda_fa_2_57_4/B sky130_fd_sc_hd__fa_1
XFILLER_39_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_423 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_34_2 dadda_fa_4_34_2/A dadda_fa_4_34_2/B dadda_fa_4_34_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_35_0/CIN dadda_fa_5_34_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_39_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_27_1 dadda_fa_4_27_1/A dadda_fa_4_27_1/B dadda_fa_4_27_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/B dadda_fa_5_27_1/B sky130_fd_sc_hd__fa_1
XFILLER_54_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ _323_/CLK _170_/D VGND VGND VPWR VPWR _170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_450 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_943 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4305 U$$4440/B1 U$$4381/A2 U$$4307/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4306/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4316 U$$4316/A U$$4366/B VGND VGND VPWR VPWR U$$4316/X sky130_fd_sc_hd__xor2_1
XU$$4327 U$$4464/A1 U$$4327/A2 U$$4466/A1 U$$4327/B2 VGND VGND VPWR VPWR U$$4328/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4338 U$$4338/A U$$4354/B VGND VGND VPWR VPWR U$$4338/X sky130_fd_sc_hd__xor2_1
XU$$4349 U$$4484/B1 U$$4349/A2 U$$4488/A1 U$$4349/B2 VGND VGND VPWR VPWR U$$4350/A
+ sky130_fd_sc_hd__a22o_1
XU$$3604 U$$4426/A1 U$$3636/A2 U$$4428/A1 U$$3636/B2 VGND VGND VPWR VPWR U$$3605/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_ha_3_16_1 U$$438/X U$$571/X VGND VGND VPWR VPWR dadda_fa_4_17_2/A dadda_ha_3_16_1/SUM
+ sky130_fd_sc_hd__ha_1
XU$$3615 U$$3615/A U$$3623/B VGND VGND VPWR VPWR U$$3615/X sky130_fd_sc_hd__xor2_1
XU$$3626 U$$4311/A1 U$$3566/X U$$4311/B1 U$$3567/X VGND VGND VPWR VPWR U$$3627/A sky130_fd_sc_hd__a22o_1
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3637 U$$3637/A U$$3637/B VGND VGND VPWR VPWR U$$3637/X sky130_fd_sc_hd__xor2_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2903 U$$26/A1 U$$2919/A2 U$$28/A1 U$$2919/B2 VGND VGND VPWR VPWR U$$2904/A sky130_fd_sc_hd__a22o_1
XU$$3648 U$$4468/B1 U$$3686/A2 U$$3648/B1 U$$3686/B2 VGND VGND VPWR VPWR U$$3649/A
+ sky130_fd_sc_hd__a22o_1
XU$$3659 U$$3659/A U$$3665/B VGND VGND VPWR VPWR U$$3659/X sky130_fd_sc_hd__xor2_1
XU$$2914 U$$2914/A U$$2996/B VGND VGND VPWR VPWR U$$2914/X sky130_fd_sc_hd__xor2_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2925 U$$3473/A1 U$$2949/A2 U$$2925/B1 U$$2949/B2 VGND VGND VPWR VPWR U$$2926/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2936 U$$2936/A U$$2968/B VGND VGND VPWR VPWR U$$2936/X sky130_fd_sc_hd__xor2_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_22_0 U$$317/X U$$450/X U$$583/X VGND VGND VPWR VPWR dadda_fa_4_23_0/B
+ dadda_fa_4_22_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_18_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2947 U$$4454/A1 U$$2949/A2 U$$2949/A1 U$$2949/B2 VGND VGND VPWR VPWR U$$2948/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 _251_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_241 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2958 U$$2958/A U$$2968/B VGND VGND VPWR VPWR U$$2958/X sky130_fd_sc_hd__xor2_1
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2969 U$$3243/A1 U$$2977/A2 U$$3108/A1 U$$2979/B2 VGND VGND VPWR VPWR U$$2970/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_252 U$$610/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_263 U$$2683/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_431 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_368_ _368_/CLK _368_/D VGND VGND VPWR VPWR _368_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_328 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4403_1778 VGND VGND VPWR VPWR U$$4403_1778/HI U$$4403/B sky130_fd_sc_hd__conb_1
X_299_ _304_/CLK _299_/D VGND VGND VPWR VPWR _299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_81_4 dadda_fa_2_81_4/A dadda_fa_2_81_4/B dadda_fa_2_81_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_1/CIN dadda_fa_3_81_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_5_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_556 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_74_3 dadda_fa_2_74_3/A dadda_fa_2_74_3/B dadda_fa_2_74_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/B dadda_fa_3_74_3/B sky130_fd_sc_hd__fa_1
XFILLER_25_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_67_2 dadda_fa_2_67_2/A dadda_fa_2_67_2/B dadda_fa_2_67_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/A dadda_fa_3_67_3/A sky130_fd_sc_hd__fa_1
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$909 final_adder.U$$138/A final_adder.U$$847/X final_adder.U$$909/B1
+ VGND VGND VPWR VPWR final_adder.U$$909/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_44_1 dadda_fa_5_44_1/A dadda_fa_5_44_1/B dadda_fa_5_44_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_45_0/B dadda_fa_7_44_0/A sky130_fd_sc_hd__fa_1
XFILLER_96_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_37_0 dadda_fa_5_37_0/A dadda_fa_5_37_0/B dadda_fa_5_37_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_38_0/A dadda_fa_6_37_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_209_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_5_111_0 dadda_fa_5_111_0/A dadda_fa_5_111_0/B dadda_fa_5_111_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_112_0/A dadda_fa_6_111_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_62_1 U$$2791/X U$$2924/X U$$3057/X VGND VGND VPWR VPWR dadda_fa_2_63_0/CIN
+ dadda_fa_2_62_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_86_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_55_0 U$$782/X U$$915/X U$$1048/X VGND VGND VPWR VPWR dadda_fa_2_56_0/B
+ dadda_fa_2_55_3/B sky130_fd_sc_hd__fa_1
XFILLER_74_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1509 U$$1644/A VGND VGND VPWR VPWR U$$1509/Y sky130_fd_sc_hd__inv_1
XFILLER_128_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_222_ _355_/CLK _222_/D VGND VGND VPWR VPWR _222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_91_3 dadda_fa_3_91_3/A dadda_fa_3_91_3/B dadda_fa_3_91_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_92_1/B dadda_fa_4_91_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_136_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_84_2 dadda_fa_3_84_2/A dadda_fa_3_84_2/B dadda_fa_3_84_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_1/A dadda_fa_4_84_2/B sky130_fd_sc_hd__fa_1
XFILLER_124_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_77_1 dadda_fa_3_77_1/A dadda_fa_3_77_1/B dadda_fa_3_77_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_0/CIN dadda_fa_4_77_2/A sky130_fd_sc_hd__fa_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_54_0 dadda_fa_6_54_0/A dadda_fa_6_54_0/B dadda_fa_6_54_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_55_0/B dadda_fa_7_54_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_88_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater409 U$$636/A2 VGND VGND VPWR VPWR U$$606/A2 sky130_fd_sc_hd__buf_4
XFILLER_78_665 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4102 U$$4102/A U$$4110/A VGND VGND VPWR VPWR U$$4102/X sky130_fd_sc_hd__xor2_1
XFILLER_38_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4113 U$$4243/B U$$4113/B VGND VGND VPWR VPWR U$$4113/X sky130_fd_sc_hd__and2_1
XU$$4124 U$$4398/A1 U$$4144/A2 U$$4400/A1 U$$4144/B2 VGND VGND VPWR VPWR U$$4125/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4135 U$$4135/A U$$4165/B VGND VGND VPWR VPWR U$$4135/X sky130_fd_sc_hd__xor2_1
XU$$3401 U$$3401/A U$$3417/B VGND VGND VPWR VPWR U$$3401/X sky130_fd_sc_hd__xor2_1
XU$$4146 U$$4146/A1 U$$4188/A2 input71/X U$$4188/B2 VGND VGND VPWR VPWR U$$4147/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3412 U$$3684/B1 U$$3416/A2 U$$3551/A1 U$$3416/B2 VGND VGND VPWR VPWR U$$3413/A
+ sky130_fd_sc_hd__a22o_1
XU$$4157 U$$4157/A U$$4243/B VGND VGND VPWR VPWR U$$4157/X sky130_fd_sc_hd__xor2_1
XU$$3423 U$$3423/A U$$3424/A VGND VGND VPWR VPWR U$$3423/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_113_2 dadda_fa_4_113_2/A dadda_fa_4_113_2/B dadda_fa_4_113_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_114_0/CIN dadda_fa_5_113_1/CIN sky130_fd_sc_hd__fa_1
XU$$4168 U$$4440/B1 U$$4176/A2 U$$4307/A1 U$$4176/B2 VGND VGND VPWR VPWR U$$4169/A
+ sky130_fd_sc_hd__a22o_1
XU$$4179 U$$4179/A U$$4189/B VGND VGND VPWR VPWR U$$4179/X sky130_fd_sc_hd__xor2_1
XU$$3434 U$$3434/A U$$3454/B VGND VGND VPWR VPWR U$$3434/X sky130_fd_sc_hd__xor2_1
XFILLER_20_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2700 U$$2700/A U$$2710/B VGND VGND VPWR VPWR U$$2700/X sky130_fd_sc_hd__xor2_1
XFILLER_206_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3445 input125/X U$$3489/A2 input126/X U$$3489/B2 VGND VGND VPWR VPWR U$$3446/A
+ sky130_fd_sc_hd__a22o_1
XU$$3456 U$$3456/A U$$3480/B VGND VGND VPWR VPWR U$$3456/X sky130_fd_sc_hd__xor2_1
XU$$2711 U$$2848/A1 U$$2711/A2 U$$2711/B1 U$$2711/B2 VGND VGND VPWR VPWR U$$2712/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_106_1 dadda_fa_4_106_1/A dadda_fa_4_106_1/B dadda_fa_4_106_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/B dadda_fa_5_106_1/B sky130_fd_sc_hd__fa_1
XU$$2722 U$$2722/A U$$2739/A VGND VGND VPWR VPWR U$$2722/X sky130_fd_sc_hd__xor2_1
XU$$3467 U$$4426/A1 U$$3503/A2 U$$4428/A1 U$$3503/B2 VGND VGND VPWR VPWR U$$3468/A
+ sky130_fd_sc_hd__a22o_1
XU$$2733 U$$3281/A1 U$$2735/A2 U$$3281/B1 U$$2735/B2 VGND VGND VPWR VPWR U$$2734/A
+ sky130_fd_sc_hd__a22o_1
XU$$3478 U$$3478/A U$$3480/B VGND VGND VPWR VPWR U$$3478/X sky130_fd_sc_hd__xor2_1
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2744 U$$2742/Y input35/X input33/X U$$2743/X U$$2740/Y VGND VGND VPWR VPWR U$$2744/X
+ sky130_fd_sc_hd__a32o_2
XU$$3489 U$$4311/A1 U$$3489/A2 U$$4311/B1 U$$3489/B2 VGND VGND VPWR VPWR U$$3490/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2755 U$$2755/A U$$2755/B VGND VGND VPWR VPWR U$$2755/X sky130_fd_sc_hd__xor2_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2766 U$$2901/B1 U$$2782/A2 U$$711/B1 U$$2782/B2 VGND VGND VPWR VPWR U$$2767/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2777 U$$2777/A U$$2869/B VGND VGND VPWR VPWR U$$2777/X sky130_fd_sc_hd__xor2_1
XU$$2788 U$$3473/A1 U$$2790/A2 U$$2925/B1 U$$2790/B2 VGND VGND VPWR VPWR U$$2789/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2799 U$$2799/A U$$2837/B VGND VGND VPWR VPWR U$$2799/X sky130_fd_sc_hd__xor2_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_127_0 dadda_fa_7_127_0/A dadda_fa_7_127_0/B dadda_fa_7_127_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_127_0/COUT _295_/D sky130_fd_sc_hd__fa_1
XFILLER_109_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_1046 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_72_0 dadda_fa_2_72_0/A dadda_fa_2_72_0/B dadda_fa_2_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_0/B dadda_fa_3_72_2/B sky130_fd_sc_hd__fa_1
XFILLER_9_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$706 final_adder.U$$706/A final_adder.U$$706/B VGND VGND VPWR VPWR
+ final_adder.U$$786/A sky130_fd_sc_hd__and2_1
Xrepeater910 input99/X VGND VGND VPWR VPWR U$$4333/B1 sky130_fd_sc_hd__buf_4
XFILLER_99_1104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$717 final_adder.U$$716/B final_adder.U$$613/X final_adder.U$$597/X
+ VGND VGND VPWR VPWR final_adder.U$$717/X sky130_fd_sc_hd__a21o_1
Xrepeater921 U$$4468/B1 VGND VGND VPWR VPWR U$$4333/A1 sky130_fd_sc_hd__buf_4
XFILLER_110_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater932 U$$3646/A1 VGND VGND VPWR VPWR U$$3644/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_57_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater943 U$$4188/B1 VGND VGND VPWR VPWR U$$80/A1 sky130_fd_sc_hd__buf_6
XFILLER_116_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater954 U$$3366/A1 VGND VGND VPWR VPWR U$$763/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_110_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater965 input92/X VGND VGND VPWR VPWR U$$3775/A1 sky130_fd_sc_hd__buf_4
Xrepeater976 U$$4456/A1 VGND VGND VPWR VPWR U$$2949/A1 sky130_fd_sc_hd__buf_4
Xrepeater987 U$$1209/B VGND VGND VPWR VPWR U$$1223/B sky130_fd_sc_hd__buf_8
XFILLER_209_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater998 U$$4178/B1 VGND VGND VPWR VPWR U$$4043/A1 sky130_fd_sc_hd__buf_4
XFILLER_37_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_595 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3990 U$$3990/A U$$4012/B VGND VGND VPWR VPWR U$$3990/X sky130_fd_sc_hd__xor2_1
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _385_/CLK sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_4_94_1 dadda_fa_4_94_1/A dadda_fa_4_94_1/B dadda_fa_4_94_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/B dadda_fa_5_94_1/B sky130_fd_sc_hd__fa_1
XFILLER_137_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_7_71_0 dadda_fa_7_71_0/A dadda_fa_7_71_0/B dadda_fa_7_71_0/CIN VGND VGND
+ VPWR VPWR _368_/D _239_/D sky130_fd_sc_hd__fa_1
XFILLER_146_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_87_0 dadda_fa_4_87_0/A dadda_fa_4_87_0/B dadda_fa_4_87_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/A dadda_fa_5_87_1/A sky130_fd_sc_hd__fa_1
Xdadda_fa_3_108_3 U$$4479/X input138/X dadda_fa_3_108_3/CIN VGND VGND VPWR VPWR dadda_fa_4_109_1/B
+ dadda_fa_4_108_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_133_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput270 output270/A VGND VGND VPWR VPWR o[111] sky130_fd_sc_hd__buf_2
XFILLER_133_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput281 output281/A VGND VGND VPWR VPWR o[121] sky130_fd_sc_hd__buf_2
Xoutput292 output292/A VGND VGND VPWR VPWR o[16] sky130_fd_sc_hd__buf_2
XFILLER_121_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3148_1744 VGND VGND VPWR VPWR U$$3148_1744/HI U$$3148/B1 sky130_fd_sc_hd__conb_1
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2007 U$$2007/A U$$2009/B VGND VGND VPWR VPWR U$$2007/X sky130_fd_sc_hd__xor2_1
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2018 U$$920/B1 U$$2052/A2 U$$787/A1 U$$2052/B2 VGND VGND VPWR VPWR U$$2019/A sky130_fd_sc_hd__a22o_1
XFILLER_210_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2029 U$$2029/A U$$2054/A VGND VGND VPWR VPWR U$$2029/X sky130_fd_sc_hd__xor2_1
XFILLER_56_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1306 U$$1306/A U$$1316/B VGND VGND VPWR VPWR U$$1306/X sky130_fd_sc_hd__xor2_1
XFILLER_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1317 U$$4055/B1 U$$1361/A2 U$$3922/A1 U$$1355/B2 VGND VGND VPWR VPWR U$$1318/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1328 U$$1328/A U$$1338/B VGND VGND VPWR VPWR U$$1328/X sky130_fd_sc_hd__xor2_1
XU$$1339 U$$2159/B1 U$$1353/A2 U$$2026/A1 U$$1238/X VGND VGND VPWR VPWR U$$1340/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_205_ _337_/CLK _205_/D VGND VGND VPWR VPWR _205_/Q sky130_fd_sc_hd__dfxtp_1
Xfinal_adder.U$$1100 final_adder.U$$178/A final_adder.U$$887/X VGND VGND VPWR VPWR
+ output358/A sky130_fd_sc_hd__xor2_1
XFILLER_128_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1111 final_adder.U$$168/B final_adder.U$$939/X VGND VGND VPWR VPWR
+ output370/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1122 final_adder.U$$156/A final_adder.U$$865/X VGND VGND VPWR VPWR
+ output382/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1133 final_adder.U$$146/B final_adder.U$$917/X VGND VGND VPWR VPWR
+ output267/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1144 final_adder.U$$134/A final_adder.U$$843/X VGND VGND VPWR VPWR
+ output280/A sky130_fd_sc_hd__xor2_1
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1000 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_960 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1022 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_504 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_930 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_51_5 dadda_fa_2_51_5/A dadda_fa_2_51_5/B dadda_fa_2_51_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_52_2/A dadda_fa_4_51_0/A sky130_fd_sc_hd__fa_1
XFILLER_93_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_955 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_44_4 dadda_fa_2_44_4/A dadda_fa_2_44_4/B dadda_fa_2_44_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_1/CIN dadda_fa_3_44_3/CIN sky130_fd_sc_hd__fa_1
XU$$3220 U$$3220/A U$$3256/B VGND VGND VPWR VPWR U$$3220/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_6_3_0 U$$13/X U$$146/X VGND VGND VPWR VPWR dadda_fa_7_4_0/B dadda_ha_6_3_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$3231 U$$3642/A1 U$$3155/X U$$3644/A1 U$$3156/X VGND VGND VPWR VPWR U$$3232/A sky130_fd_sc_hd__a22o_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$13 _309_/Q _181_/Q VGND VGND VPWR VPWR final_adder.U$$243/B1 final_adder.U$$242/B
+ sky130_fd_sc_hd__ha_1
XU$$3242 U$$3242/A U$$3242/B VGND VGND VPWR VPWR U$$3242/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$24 _320_/Q _192_/Q VGND VGND VPWR VPWR final_adder.U$$231/A2 final_adder.U$$230/A
+ sky130_fd_sc_hd__ha_1
XU$$3253 U$$650/A1 U$$3255/A2 U$$789/A1 U$$3255/B2 VGND VGND VPWR VPWR U$$3254/A sky130_fd_sc_hd__a22o_1
XFILLER_19_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$35 _331_/Q _203_/Q VGND VGND VPWR VPWR final_adder.U$$221/B1 final_adder.U$$220/B
+ sky130_fd_sc_hd__ha_1
XU$$3264 U$$3264/A U$$3264/B VGND VGND VPWR VPWR U$$3264/X sky130_fd_sc_hd__xor2_1
XFILLER_47_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_37_3 U$$1943/X U$$2076/X U$$2209/X VGND VGND VPWR VPWR dadda_fa_3_38_1/B
+ dadda_fa_3_37_3/B sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$46 _342_/Q _214_/Q VGND VGND VPWR VPWR final_adder.U$$979/B1 final_adder.U$$208/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3275 U$$3684/B1 U$$3277/A2 U$$3551/A1 U$$3277/B2 VGND VGND VPWR VPWR U$$3276/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$57 _353_/Q _225_/Q VGND VGND VPWR VPWR final_adder.U$$199/B1 final_adder.U$$198/B
+ sky130_fd_sc_hd__ha_1
XU$$2530 U$$3352/A1 U$$2558/A2 U$$3078/B1 U$$2558/B2 VGND VGND VPWR VPWR U$$2531/A
+ sky130_fd_sc_hd__a22o_1
XU$$3286 U$$3286/A U$$3286/B VGND VGND VPWR VPWR U$$3286/X sky130_fd_sc_hd__xor2_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2541 U$$2541/A U$$2569/B VGND VGND VPWR VPWR U$$2541/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$68 _364_/Q _236_/Q VGND VGND VPWR VPWR final_adder.U$$957/B1 final_adder.U$$186/A
+ sky130_fd_sc_hd__ha_1
XU$$2552 U$$3922/A1 U$$2600/A2 U$$3922/B1 U$$2600/B2 VGND VGND VPWR VPWR U$$2553/A
+ sky130_fd_sc_hd__a22o_1
XU$$3297 U$$3297/A U$$3321/B VGND VGND VPWR VPWR U$$3297/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$79 _375_/Q _247_/Q VGND VGND VPWR VPWR final_adder.U$$177/B1 final_adder.U$$176/B
+ sky130_fd_sc_hd__ha_1
XFILLER_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2563 U$$2563/A U$$2603/A VGND VGND VPWR VPWR U$$2563/X sky130_fd_sc_hd__xor2_1
XU$$2574 U$$2709/B1 U$$2576/A2 U$$2711/B1 U$$2576/B2 VGND VGND VPWR VPWR U$$2575/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1840 U$$1840/A U$$1840/B VGND VGND VPWR VPWR U$$1840/X sky130_fd_sc_hd__xor2_1
XU$$2585 U$$2585/A U$$2602/A VGND VGND VPWR VPWR U$$2585/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2596 U$$3281/A1 U$$2596/A2 U$$3281/B1 U$$2596/B2 VGND VGND VPWR VPWR U$$2597/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1851 U$$616/B1 U$$1879/A2 U$$2949/A1 U$$1879/B2 VGND VGND VPWR VPWR U$$1852/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1862 U$$1862/A U$$1870/B VGND VGND VPWR VPWR U$$1862/X sky130_fd_sc_hd__xor2_1
XFILLER_107_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1873 U$$2967/B1 U$$1877/A2 U$$94/A1 U$$1877/B2 VGND VGND VPWR VPWR U$$1874/A sky130_fd_sc_hd__a22o_1
XFILLER_21_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1884 U$$1884/A U$$1914/B VGND VGND VPWR VPWR U$$1884/X sky130_fd_sc_hd__xor2_1
XFILLER_166_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1895 U$$2032/A1 U$$1915/A2 U$$2582/A1 U$$1915/B2 VGND VGND VPWR VPWR U$$1896/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_478 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$503 final_adder.U$$498/A final_adder.U$$381/X final_adder.U$$377/X
+ VGND VGND VPWR VPWR final_adder.U$$503/X sky130_fd_sc_hd__a21o_2
XTAP_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$514 final_adder.U$$522/B final_adder.U$$514/B VGND VGND VPWR VPWR
+ final_adder.U$$634/B sky130_fd_sc_hd__and2_1
XFILLER_97_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$525 final_adder.U$$524/B final_adder.U$$409/X final_adder.U$$401/X
+ VGND VGND VPWR VPWR final_adder.U$$525/X sky130_fd_sc_hd__a21o_1
XFILLER_9_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_635 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$536 final_adder.U$$544/B final_adder.U$$536/B VGND VGND VPWR VPWR
+ final_adder.U$$656/B sky130_fd_sc_hd__and2_1
XTAP_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater740 U$$3293/X VGND VGND VPWR VPWR U$$3374/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$547 final_adder.U$$546/B final_adder.U$$431/X final_adder.U$$423/X
+ VGND VGND VPWR VPWR final_adder.U$$547/X sky130_fd_sc_hd__a21o_1
XTAP_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater751 U$$3098/B2 VGND VGND VPWR VPWR U$$3108/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$558 final_adder.U$$566/B final_adder.U$$558/B VGND VGND VPWR VPWR
+ final_adder.U$$678/B sky130_fd_sc_hd__and2_1
XTAP_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater762 U$$2967/B2 VGND VGND VPWR VPWR U$$2949/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$569 final_adder.U$$568/B final_adder.U$$453/X final_adder.U$$445/X
+ VGND VGND VPWR VPWR final_adder.U$$569/X sky130_fd_sc_hd__a21o_1
XU$$408 U$$817/B1 U$$278/X U$$408/B1 U$$279/X VGND VGND VPWR VPWR U$$409/A sky130_fd_sc_hd__a22o_1
Xrepeater773 U$$279/X VGND VGND VPWR VPWR U$$396/B2 sky130_fd_sc_hd__buf_4
XU$$419 U$$8/A1 U$$437/A2 U$$8/B1 U$$437/B2 VGND VGND VPWR VPWR U$$420/A sky130_fd_sc_hd__a22o_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater784 U$$2683/B2 VGND VGND VPWR VPWR U$$2653/B2 sky130_fd_sc_hd__buf_4
Xrepeater795 U$$2542/B2 VGND VGND VPWR VPWR U$$2524/B2 sky130_fd_sc_hd__buf_6
XFILLER_38_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2052_1726 VGND VGND VPWR VPWR U$$2052_1726/HI U$$2052/B1 sky130_fd_sc_hd__conb_1
XFILLER_38_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1308 U$$3425/A VGND VGND VPWR VPWR U$$3389/B sky130_fd_sc_hd__buf_6
XFILLER_119_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_3_113_1 U$$3824/X U$$3957/X U$$4090/X VGND VGND VPWR VPWR dadda_fa_4_114_2/A
+ dadda_fa_4_113_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater1319 U$$3288/A VGND VGND VPWR VPWR U$$3256/B sky130_fd_sc_hd__buf_6
XFILLER_114_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_106_0 U$$3544/X U$$3677/X U$$3810/X VGND VGND VPWR VPWR dadda_fa_4_107_0/B
+ dadda_fa_4_106_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_109_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_54_3 dadda_fa_3_54_3/A dadda_fa_3_54_3/B dadda_fa_3_54_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_55_1/B dadda_fa_4_54_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_94_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_47_2 dadda_fa_3_47_2/A dadda_fa_3_47_2/B dadda_fa_3_47_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_1/A dadda_fa_4_47_2/B sky130_fd_sc_hd__fa_1
XFILLER_29_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_80_0_1852 VGND VGND VPWR VPWR dadda_fa_1_80_0/A dadda_fa_1_80_0_1852/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_63_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$920 U$$920/A1 U$$950/A2 U$$920/B1 U$$950/B2 VGND VGND VPWR VPWR U$$921/A sky130_fd_sc_hd__a22o_1
XU$$931 U$$931/A U$$945/B VGND VGND VPWR VPWR U$$931/X sky130_fd_sc_hd__xor2_1
XU$$942 U$$942/A1 U$$950/A2 U$$944/A1 U$$950/B2 VGND VGND VPWR VPWR U$$943/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_6_17_0 dadda_fa_6_17_0/A dadda_fa_6_17_0/B dadda_fa_6_17_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_18_0/B dadda_fa_7_17_0/CIN sky130_fd_sc_hd__fa_1
XU$$953 U$$953/A U$$958/A VGND VGND VPWR VPWR U$$953/X sky130_fd_sc_hd__xor2_1
XU$$1103 U$$1103/A U$$1139/B VGND VGND VPWR VPWR U$$1103/X sky130_fd_sc_hd__xor2_1
XFILLER_141_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$964 U$$962/B input5/X input6/X U$$959/Y VGND VGND VPWR VPWR U$$964/X sky130_fd_sc_hd__a22o_2
XU$$1114 U$$3032/A1 U$$1138/A2 U$$979/A1 U$$1138/B2 VGND VGND VPWR VPWR U$$1115/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$975 U$$975/A1 U$$979/A2 U$$18/A1 U$$979/B2 VGND VGND VPWR VPWR U$$976/A sky130_fd_sc_hd__a22o_1
XU$$1125 U$$1125/A U$$1137/B VGND VGND VPWR VPWR U$$1125/X sky130_fd_sc_hd__xor2_1
XU$$986 U$$986/A U$$996/B VGND VGND VPWR VPWR U$$986/X sky130_fd_sc_hd__xor2_1
XFILLER_44_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$997 U$$997/A1 U$$997/A2 U$$997/B1 U$$997/B2 VGND VGND VPWR VPWR U$$998/A sky130_fd_sc_hd__a22o_1
XU$$1136 U$$999/A1 U$$1136/A2 U$$42/A1 U$$1136/B2 VGND VGND VPWR VPWR U$$1137/A sky130_fd_sc_hd__a22o_1
XU$$1147 U$$1147/A U$$1187/B VGND VGND VPWR VPWR U$$1147/X sky130_fd_sc_hd__xor2_1
XU$$1158 U$$62/A1 U$$1162/A2 U$$62/B1 U$$1162/B2 VGND VGND VPWR VPWR U$$1159/A sky130_fd_sc_hd__a22o_1
XU$$1169 U$$1169/A U$$1175/B VGND VGND VPWR VPWR U$$1169/X sky130_fd_sc_hd__xor2_1
XFILLER_70_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_42_1 U$$2352/X U$$2485/X U$$2618/X VGND VGND VPWR VPWR dadda_fa_3_43_0/CIN
+ dadda_fa_3_42_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_38_167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3050 U$$4144/B1 U$$3082/A2 U$$4011/A1 U$$3082/B2 VGND VGND VPWR VPWR U$$3051/A
+ sky130_fd_sc_hd__a22o_1
XU$$3061 U$$3061/A U$$3077/B VGND VGND VPWR VPWR U$$3061/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_0 U$$343/X U$$476/X U$$609/X VGND VGND VPWR VPWR dadda_fa_3_36_0/B
+ dadda_fa_3_35_2/B sky130_fd_sc_hd__fa_1
XU$$3072 U$$4442/A1 U$$3098/A2 U$$4442/B1 U$$3098/B2 VGND VGND VPWR VPWR U$$3073/A
+ sky130_fd_sc_hd__a22o_1
XU$$3083 U$$3083/A U$$3083/B VGND VGND VPWR VPWR U$$3083/X sky130_fd_sc_hd__xor2_1
XFILLER_34_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3094 U$$3642/A1 U$$3018/X U$$3644/A1 U$$3019/X VGND VGND VPWR VPWR U$$3095/A sky130_fd_sc_hd__a22o_1
XU$$2360 U$$2360/A U$$2360/B VGND VGND VPWR VPWR U$$2360/X sky130_fd_sc_hd__xor2_1
XU$$2371 U$$4013/B1 U$$2463/A2 U$$4015/B1 U$$2463/B2 VGND VGND VPWR VPWR U$$2372/A
+ sky130_fd_sc_hd__a22o_1
XU$$2382 U$$2382/A U$$2465/A VGND VGND VPWR VPWR U$$2382/X sky130_fd_sc_hd__xor2_1
XFILLER_62_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2393 U$$62/B1 U$$2403/A2 U$$888/A1 U$$2403/B2 VGND VGND VPWR VPWR U$$2394/A sky130_fd_sc_hd__a22o_1
XFILLER_195_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1670 U$$983/B1 U$$1706/A2 U$$850/A1 U$$1706/B2 VGND VGND VPWR VPWR U$$1671/A sky130_fd_sc_hd__a22o_1
XFILLER_194_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1681 U$$1681/A U$$1689/B VGND VGND VPWR VPWR U$$1681/X sky130_fd_sc_hd__xor2_1
XFILLER_10_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1692 U$$3473/A1 U$$1746/A2 U$$2925/B1 U$$1746/B2 VGND VGND VPWR VPWR U$$1693/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_721 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_554 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_87_3 U$$2841/X U$$2974/X U$$3107/X VGND VGND VPWR VPWR dadda_fa_2_88_4/A
+ dadda_fa_2_87_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_1_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_64_2 dadda_fa_4_64_2/A dadda_fa_4_64_2/B dadda_fa_4_64_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_65_0/CIN dadda_fa_5_64_1/CIN sky130_fd_sc_hd__fa_1
XTAP_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_57_1 dadda_fa_4_57_1/A dadda_fa_4_57_1/B dadda_fa_4_57_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/B dadda_fa_5_57_1/B sky130_fd_sc_hd__fa_1
XFILLER_39_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfinal_adder.U$$300 final_adder.U$$302/B final_adder.U$$300/B VGND VGND VPWR VPWR
+ final_adder.U$$426/B sky130_fd_sc_hd__and2_1
XTAP_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$311 final_adder.U$$310/B final_adder.U$$185/X final_adder.U$$183/X
+ VGND VGND VPWR VPWR final_adder.U$$311/X sky130_fd_sc_hd__a21o_1
XTAP_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_34_0 dadda_fa_7_34_0/A dadda_fa_7_34_0/B dadda_fa_7_34_0/CIN VGND VGND
+ VPWR VPWR _331_/D _202_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$322 final_adder.U$$324/B final_adder.U$$322/B VGND VGND VPWR VPWR
+ final_adder.U$$448/B sky130_fd_sc_hd__and2_1
XTAP_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$333 final_adder.U$$332/B final_adder.U$$207/X final_adder.U$$205/X
+ VGND VGND VPWR VPWR final_adder.U$$333/X sky130_fd_sc_hd__a21o_1
XTAP_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$344 final_adder.U$$346/B final_adder.U$$344/B VGND VGND VPWR VPWR
+ final_adder.U$$470/B sky130_fd_sc_hd__and2_1
XTAP_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$355 final_adder.U$$354/B final_adder.U$$229/X final_adder.U$$227/X
+ VGND VGND VPWR VPWR final_adder.U$$355/X sky130_fd_sc_hd__a21o_1
XTAP_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_999 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$366 final_adder.U$$368/B final_adder.U$$366/B VGND VGND VPWR VPWR
+ final_adder.U$$492/B sky130_fd_sc_hd__and2_1
XTAP_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater570 U$$2149/A2 VGND VGND VPWR VPWR U$$2099/A2 sky130_fd_sc_hd__buf_4
XFILLER_85_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$205 U$$68/A1 U$$209/A2 U$$70/A1 U$$209/B2 VGND VGND VPWR VPWR U$$206/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$377 final_adder.U$$376/B final_adder.U$$251/X final_adder.U$$249/X
+ VGND VGND VPWR VPWR final_adder.U$$377/X sky130_fd_sc_hd__a21o_1
XTAP_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater581 U$$2040/A2 VGND VGND VPWR VPWR U$$1960/A2 sky130_fd_sc_hd__buf_4
XU$$216 U$$216/A U$$218/B VGND VGND VPWR VPWR U$$216/X sky130_fd_sc_hd__xor2_1
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$388 final_adder.U$$392/B final_adder.U$$388/B VGND VGND VPWR VPWR
+ final_adder.U$$512/B sky130_fd_sc_hd__and2_2
XTAP_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater592 U$$1736/A2 VGND VGND VPWR VPWR U$$1688/A2 sky130_fd_sc_hd__buf_4
XU$$227 U$$90/A1 U$$263/A2 U$$92/A1 U$$231/B2 VGND VGND VPWR VPWR U$$228/A sky130_fd_sc_hd__a22o_1
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$399 final_adder.U$$398/B final_adder.U$$277/X final_adder.U$$273/X
+ VGND VGND VPWR VPWR final_adder.U$$399/X sky130_fd_sc_hd__a21o_1
XU$$238 U$$238/A U$$244/B VGND VGND VPWR VPWR U$$238/X sky130_fd_sc_hd__xor2_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$249 U$$384/B1 U$$257/A2 U$$251/A1 U$$257/B2 VGND VGND VPWR VPWR U$$250/A sky130_fd_sc_hd__a22o_1
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_304 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1051 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1105 input76/X VGND VGND VPWR VPWR U$$4394/A1 sky130_fd_sc_hd__buf_4
XFILLER_154_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1116 U$$3878/B1 VGND VGND VPWR VPWR U$$3058/A1 sky130_fd_sc_hd__buf_6
Xrepeater1127 U$$4426/A1 VGND VGND VPWR VPWR U$$3876/B1 sky130_fd_sc_hd__buf_8
Xrepeater1138 U$$312/A1 VGND VGND VPWR VPWR U$$38/A1 sky130_fd_sc_hd__buf_4
XFILLER_153_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1149 U$$4144/B1 VGND VGND VPWR VPWR U$$995/A1 sky130_fd_sc_hd__buf_6
XFILLER_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_1134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_0_75_1 U$$1221/X U$$1354/X U$$1487/X VGND VGND VPWR VPWR dadda_fa_1_76_8/B
+ dadda_fa_2_75_0/A sky130_fd_sc_hd__fa_2
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_52_0 dadda_fa_3_52_0/A dadda_fa_3_52_0/B dadda_fa_3_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_0/B dadda_fa_4_52_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_68_0 dadda_fa_0_68_0/A U$$409/X U$$542/X VGND VGND VPWR VPWR dadda_fa_1_69_5/CIN
+ dadda_fa_1_68_7/B sky130_fd_sc_hd__fa_1
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$750 U$$750/A U$$750/B VGND VGND VPWR VPWR U$$750/X sky130_fd_sc_hd__xor2_1
XFILLER_95_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$761 U$$896/B1 U$$805/A2 U$$763/A1 U$$805/B2 VGND VGND VPWR VPWR U$$762/A sky130_fd_sc_hd__a22o_1
XFILLER_205_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$772 U$$772/A U$$794/B VGND VGND VPWR VPWR U$$772/X sky130_fd_sc_hd__xor2_1
XU$$783 U$$783/A1 U$$783/A2 U$$783/B1 U$$783/B2 VGND VGND VPWR VPWR U$$784/A sky130_fd_sc_hd__a22o_1
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$794 U$$794/A U$$794/B VGND VGND VPWR VPWR U$$794/X sky130_fd_sc_hd__xor2_1
XFILLER_177_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_816 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_0 ANTENNA_0/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_2_97_2 U$$3127/X U$$3260/X U$$3393/X VGND VGND VPWR VPWR dadda_fa_3_98_1/A
+ dadda_fa_3_97_3/A sky130_fd_sc_hd__fa_1
XFILLER_104_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1650 U$$789/A1 VGND VGND VPWR VPWR U$$3116/B1 sky130_fd_sc_hd__buf_8
Xdadda_fa_5_74_1 dadda_fa_5_74_1/A dadda_fa_5_74_1/B dadda_fa_5_74_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_75_0/B dadda_fa_7_74_0/A sky130_fd_sc_hd__fa_1
Xrepeater1661 U$$4484/A1 VGND VGND VPWR VPWR U$$4210/A1 sky130_fd_sc_hd__buf_4
XFILLER_132_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1672 U$$2016/A1 VGND VGND VPWR VPWR U$$2975/A1 sky130_fd_sc_hd__buf_6
Xrepeater1683 input103/X VGND VGND VPWR VPWR U$$3245/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_141_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1694 U$$914/A1 VGND VGND VPWR VPWR U$$640/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_67_0 dadda_fa_5_67_0/A dadda_fa_5_67_0/B dadda_fa_5_67_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_68_0/A dadda_fa_6_67_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_63_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_66_8 dadda_fa_1_66_8/A dadda_fa_1_66_8/B dadda_fa_1_66_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_67_3/A dadda_fa_3_66_0/A sky130_fd_sc_hd__fa_2
XFILLER_86_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_59_7 dadda_fa_1_59_7/A dadda_fa_1_59_7/B dadda_fa_1_59_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_60_2/CIN dadda_fa_2_59_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_132_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_6_6_0 input223/X dadda_fa_6_6_0/B dadda_fa_6_6_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_7_7_0/B dadda_fa_7_6_0/CIN sky130_fd_sc_hd__fa_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2190 U$$2190/A U$$2191/A VGND VGND VPWR VPWR U$$2190/X sky130_fd_sc_hd__xor2_1
XFILLER_35_1208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_92_1 U$$2319/X U$$2452/X U$$2585/X VGND VGND VPWR VPWR dadda_fa_2_93_5/A
+ dadda_fa_2_92_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_0 U$$1506/Y U$$1640/X U$$1773/X VGND VGND VPWR VPWR dadda_fa_2_86_2/B
+ dadda_fa_2_85_4/B sky130_fd_sc_hd__fa_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4509 U$$4509/A U$$4509/B VGND VGND VPWR VPWR U$$4509/X sky130_fd_sc_hd__xor2_1
XTAP_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$130 final_adder.U$$130/A final_adder.U$$130/B VGND VGND VPWR VPWR
+ final_adder.U$$258/B sky130_fd_sc_hd__and2_1
XU$$3808 U$$3808/A U$$3826/B VGND VGND VPWR VPWR U$$3808/X sky130_fd_sc_hd__xor2_1
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$141 final_adder.U$$140/B final_adder.U$$911/B1 final_adder.U$$141/B1
+ VGND VGND VPWR VPWR final_adder.U$$141/X sky130_fd_sc_hd__a21o_1
XU$$3819 input116/X U$$3819/A2 input117/X U$$3819/B2 VGND VGND VPWR VPWR U$$3820/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$152 final_adder.U$$152/A final_adder.U$$152/B VGND VGND VPWR VPWR
+ final_adder.U$$280/B sky130_fd_sc_hd__and2_1
XTAP_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$163 final_adder.U$$162/B final_adder.U$$933/B1 final_adder.U$$163/B1
+ VGND VGND VPWR VPWR final_adder.U$$163/X sky130_fd_sc_hd__a21o_1
XTAP_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$174 final_adder.U$$174/A final_adder.U$$174/B VGND VGND VPWR VPWR
+ final_adder.U$$302/B sky130_fd_sc_hd__and2_1
XTAP_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$185 final_adder.U$$184/B final_adder.U$$955/B1 final_adder.U$$185/B1
+ VGND VGND VPWR VPWR final_adder.U$$185/X sky130_fd_sc_hd__a21o_1
XTAP_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$196 final_adder.U$$196/A final_adder.U$$196/B VGND VGND VPWR VPWR
+ final_adder.U$$324/B sky130_fd_sc_hd__and2_1
XTAP_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_ha_5_126_0 dadda_ha_5_126_0/A U$$4382/X VGND VGND VPWR VPWR dadda_fa_7_127_0/A
+ dadda_fa_7_126_0/A sky130_fd_sc_hd__ha_1
XFILLER_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_52_clk _239_/CLK VGND VGND VPWR VPWR _373_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_158_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_384_ _384_/CLK _384_/D VGND VGND VPWR VPWR _384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_899 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_6_84_0 dadda_fa_6_84_0/A dadda_fa_6_84_0/B dadda_fa_6_84_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_85_0/B dadda_fa_7_84_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_495 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$134_1714 VGND VGND VPWR VPWR U$$134_1714/HI U$$134/B1 sky130_fd_sc_hd__conb_1
XFILLER_23_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput170 c[21] VGND VGND VPWR VPWR input170/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput181 c[31] VGND VGND VPWR VPWR input181/X sky130_fd_sc_hd__buf_2
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput192 c[41] VGND VGND VPWR VPWR input192/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$580 U$$717/A1 U$$606/A2 U$$34/A1 U$$606/B2 VGND VGND VPWR VPWR U$$581/A sky130_fd_sc_hd__a22o_1
XFILLER_211_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$591 U$$591/A U$$625/B VGND VGND VPWR VPWR U$$591/X sky130_fd_sc_hd__xor2_1
XFILLER_51_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_43_clk _385_/CLK VGND VGND VPWR VPWR _382_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1480 input126/X VGND VGND VPWR VPWR U$$4406/A1 sky130_fd_sc_hd__buf_6
Xrepeater1491 U$$3283/B1 VGND VGND VPWR VPWR U$$956/A1 sky130_fd_sc_hd__buf_4
XFILLER_87_803 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3285_1746 VGND VGND VPWR VPWR U$$3285_1746/HI U$$3285/B1 sky130_fd_sc_hd__conb_1
XFILLER_8_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_71_6 input225/X dadda_fa_1_71_6/B dadda_fa_1_71_6/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_72_2/B dadda_fa_2_71_5/B sky130_fd_sc_hd__fa_1
XFILLER_99_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_64_5 input217/X dadda_fa_1_64_5/B dadda_fa_1_64_5/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_65_2/A dadda_fa_2_64_5/A sky130_fd_sc_hd__fa_1
XFILLER_87_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_1_57_4 U$$2781/X U$$2914/X U$$3047/X VGND VGND VPWR VPWR dadda_fa_2_58_1/CIN
+ dadda_fa_2_57_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_27_2 dadda_fa_4_27_2/A dadda_fa_4_27_2/B dadda_fa_4_27_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_28_0/CIN dadda_fa_5_27_1/CIN sky130_fd_sc_hd__fa_1
XU$$4461_1807 VGND VGND VPWR VPWR U$$4461_1807/HI U$$4461/B sky130_fd_sc_hd__conb_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1025 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_73 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_462 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4306 U$$4306/A U$$4384/A VGND VGND VPWR VPWR U$$4306/X sky130_fd_sc_hd__xor2_1
XFILLER_120_966 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4317 U$$4454/A1 U$$4327/A2 U$$4456/A1 U$$4327/B2 VGND VGND VPWR VPWR U$$4318/A
+ sky130_fd_sc_hd__a22o_1
XU$$4328 U$$4328/A U$$4330/B VGND VGND VPWR VPWR U$$4328/X sky130_fd_sc_hd__xor2_1
XU$$4339 input101/X U$$4349/A2 U$$4478/A1 U$$4349/B2 VGND VGND VPWR VPWR U$$4340/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_936 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3605 U$$3605/A U$$3637/B VGND VGND VPWR VPWR U$$3605/X sky130_fd_sc_hd__xor2_1
XU$$3616 input80/X U$$3660/A2 input81/X U$$3660/B2 VGND VGND VPWR VPWR U$$3617/A sky130_fd_sc_hd__a22o_1
XU$$3627 U$$3627/A input49/X VGND VGND VPWR VPWR U$$3627/X sky130_fd_sc_hd__xor2_1
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3638 U$$3775/A1 U$$3566/X U$$3775/B1 U$$3567/X VGND VGND VPWR VPWR U$$3639/A sky130_fd_sc_hd__a22o_1
XFILLER_46_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2904 U$$2904/A U$$2920/B VGND VGND VPWR VPWR U$$2904/X sky130_fd_sc_hd__xor2_1
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3649 U$$3649/A U$$3697/B VGND VGND VPWR VPWR U$$3649/X sky130_fd_sc_hd__xor2_1
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2915 U$$4011/A1 U$$2919/A2 U$$38/B1 U$$2919/B2 VGND VGND VPWR VPWR U$$2916/A sky130_fd_sc_hd__a22o_1
XU$$2926 U$$2926/A U$$2950/B VGND VGND VPWR VPWR U$$2926/X sky130_fd_sc_hd__xor2_1
XFILLER_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_220 _213_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2937 U$$4442/B1 U$$2967/A2 U$$3211/B1 U$$2967/B2 VGND VGND VPWR VPWR U$$2938/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2948 U$$2948/A U$$2950/B VGND VGND VPWR VPWR U$$2948/X sky130_fd_sc_hd__xor2_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2959 U$$3644/A1 U$$2985/A2 U$$3644/B1 U$$2985/B2 VGND VGND VPWR VPWR U$$2960/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_22_1 U$$716/X U$$849/X U$$982/X VGND VGND VPWR VPWR dadda_fa_4_23_0/CIN
+ dadda_fa_4_22_2/A sky130_fd_sc_hd__fa_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_242 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 input109/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_264 U$$2302/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk _380_/CLK VGND VGND VPWR VPWR _384_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_367_ _367_/CLK _367_/D VGND VGND VPWR VPWR _367_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_298_ _323_/CLK _298_/D VGND VGND VPWR VPWR _298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_81_5 dadda_fa_2_81_5/A dadda_fa_2_81_5/B dadda_fa_2_81_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_82_2/A dadda_fa_4_81_0/A sky130_fd_sc_hd__fa_2
XFILLER_114_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_74_4 dadda_fa_2_74_4/A dadda_fa_2_74_4/B dadda_fa_2_74_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_1/CIN dadda_fa_3_74_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_67_3 dadda_fa_2_67_3/A dadda_fa_2_67_3/B dadda_fa_2_67_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/B dadda_fa_3_67_3/B sky130_fd_sc_hd__fa_1
XFILLER_110_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_37_1 dadda_fa_5_37_1/A dadda_fa_5_37_1/B dadda_fa_5_37_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_38_0/B dadda_fa_7_37_0/A sky130_fd_sc_hd__fa_1
XFILLER_83_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_209_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk _227_/CLK VGND VGND VPWR VPWR _357_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_111_1 dadda_fa_5_111_1/A dadda_fa_5_111_1/B dadda_fa_5_111_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_112_0/B dadda_fa_7_111_0/A sky130_fd_sc_hd__fa_1
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_104_0 dadda_fa_5_104_0/A dadda_fa_5_104_0/B dadda_fa_5_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_105_0/A dadda_fa_6_104_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_1096 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4419_1786 VGND VGND VPWR VPWR U$$4419_1786/HI U$$4419/B sky130_fd_sc_hd__conb_1
XFILLER_161_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_62_2 U$$3190/X U$$3323/X U$$3456/X VGND VGND VPWR VPWR dadda_fa_2_63_1/A
+ dadda_fa_2_62_4/A sky130_fd_sc_hd__fa_1
XFILLER_101_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_55_1 U$$1181/X U$$1314/X U$$1447/X VGND VGND VPWR VPWR dadda_fa_2_56_0/CIN
+ dadda_fa_2_55_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_170_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_32_0 dadda_fa_4_32_0/A dadda_fa_4_32_0/B dadda_fa_4_32_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/A dadda_fa_5_32_1/A sky130_fd_sc_hd__fa_1
XFILLER_132_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_48_0 U$$103/X U$$236/X U$$369/X VGND VGND VPWR VPWR dadda_fa_2_49_1/A
+ dadda_fa_2_48_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_16_928 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_221_ _351_/CLK _221_/D VGND VGND VPWR VPWR _221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_84_3 dadda_fa_3_84_3/A dadda_fa_3_84_3/B dadda_fa_3_84_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_85_1/B dadda_fa_4_84_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_163_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_77_2 dadda_fa_3_77_2/A dadda_fa_3_77_2/B dadda_fa_3_77_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_1/A dadda_fa_4_77_2/B sky130_fd_sc_hd__fa_1
XFILLER_105_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_47_0 dadda_fa_6_47_0/A dadda_fa_6_47_0/B dadda_fa_6_47_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_48_0/B dadda_fa_7_47_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_78_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4103 U$$4375/B1 U$$4103/A2 U$$4103/B1 U$$4103/B2 VGND VGND VPWR VPWR U$$4104/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4114 U$$4112/Y input57/X input55/X U$$4113/X U$$4110/Y VGND VGND VPWR VPWR U$$4114/X
+ sky130_fd_sc_hd__a32o_2
XU$$4125 U$$4125/A U$$4145/B VGND VGND VPWR VPWR U$$4125/X sky130_fd_sc_hd__xor2_1
XFILLER_66_839 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4136 U$$4273/A1 U$$4164/A2 U$$4273/B1 U$$4164/B2 VGND VGND VPWR VPWR U$$4137/A
+ sky130_fd_sc_hd__a22o_1
XU$$3402 input113/X U$$3422/A2 input114/X U$$3422/B2 VGND VGND VPWR VPWR U$$3403/A
+ sky130_fd_sc_hd__a22o_1
XU$$4147 U$$4147/A U$$4189/B VGND VGND VPWR VPWR U$$4147/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3413 U$$3413/A U$$3417/B VGND VGND VPWR VPWR U$$3413/X sky130_fd_sc_hd__xor2_1
XFILLER_24_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4158 U$$4293/B1 U$$4164/A2 input78/X U$$4164/B2 VGND VGND VPWR VPWR U$$4159/A
+ sky130_fd_sc_hd__a22o_1
XU$$3424 U$$3424/A VGND VGND VPWR VPWR U$$3424/Y sky130_fd_sc_hd__inv_1
XU$$4169 U$$4169/A U$$4246/A VGND VGND VPWR VPWR U$$4169/X sky130_fd_sc_hd__xor2_1
XU$$3435 U$$832/A1 U$$3527/A2 U$$3846/B1 U$$3527/B2 VGND VGND VPWR VPWR U$$3436/A
+ sky130_fd_sc_hd__a22o_1
XU$$3446 U$$3446/A U$$3490/B VGND VGND VPWR VPWR U$$3446/X sky130_fd_sc_hd__xor2_1
XU$$2701 U$$2975/A1 U$$2711/A2 U$$2701/B1 U$$2711/B2 VGND VGND VPWR VPWR U$$2702/A
+ sky130_fd_sc_hd__a22o_1
XU$$3457 U$$3594/A1 U$$3479/A2 U$$4005/B1 U$$3479/B2 VGND VGND VPWR VPWR U$$3458/A
+ sky130_fd_sc_hd__a22o_1
XU$$2712 U$$2712/A input33/X VGND VGND VPWR VPWR U$$2712/X sky130_fd_sc_hd__xor2_1
XFILLER_92_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_106_2 dadda_fa_4_106_2/A dadda_fa_4_106_2/B dadda_fa_4_106_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_107_0/CIN dadda_fa_5_106_1/CIN sky130_fd_sc_hd__fa_1
XU$$2723 U$$118/B1 U$$2735/A2 U$$122/A1 U$$2735/B2 VGND VGND VPWR VPWR U$$2724/A sky130_fd_sc_hd__a22o_1
XFILLER_111_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3468 U$$3468/A U$$3504/B VGND VGND VPWR VPWR U$$3468/X sky130_fd_sc_hd__xor2_1
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2734 U$$2734/A U$$2736/B VGND VGND VPWR VPWR U$$2734/X sky130_fd_sc_hd__xor2_1
XU$$3479 U$$4027/A1 U$$3479/A2 U$$741/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3480/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2745 U$$2743/B input33/X input35/X U$$2740/Y VGND VGND VPWR VPWR U$$2745/X sky130_fd_sc_hd__a22o_2
XFILLER_209_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2756 U$$3987/B1 U$$2790/A2 U$$3852/B1 U$$2790/B2 VGND VGND VPWR VPWR U$$2757/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2767 U$$2767/A U$$2783/B VGND VGND VPWR VPWR U$$2767/X sky130_fd_sc_hd__xor2_1
XFILLER_2_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2778 U$$312/A1 U$$2782/A2 U$$38/B1 U$$2782/B2 VGND VGND VPWR VPWR U$$2779/A sky130_fd_sc_hd__a22o_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2789 U$$2789/A U$$2797/B VGND VGND VPWR VPWR U$$2789/X sky130_fd_sc_hd__xor2_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_419_ _419_/CLK _419_/D VGND VGND VPWR VPWR _419_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_811 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _326_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_72_1 dadda_fa_2_72_1/A dadda_fa_2_72_1/B dadda_fa_2_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_0/CIN dadda_fa_3_72_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_65_0 dadda_fa_2_65_0/A dadda_fa_2_65_0/B dadda_fa_2_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_0/B dadda_fa_3_65_2/B sky130_fd_sc_hd__fa_1
Xrepeater900 U$$4498/B2 VGND VGND VPWR VPWR U$$4494/B2 sky130_fd_sc_hd__buf_4
XFILLER_57_806 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$707 final_adder.U$$706/B final_adder.U$$603/X final_adder.U$$587/X
+ VGND VGND VPWR VPWR final_adder.U$$707/X sky130_fd_sc_hd__a21o_1
Xrepeater911 U$$836/A1 VGND VGND VPWR VPWR U$$14/A1 sky130_fd_sc_hd__buf_6
XFILLER_111_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$718 final_adder.U$$718/A final_adder.U$$718/B VGND VGND VPWR VPWR
+ final_adder.U$$798/A sky130_fd_sc_hd__and2_1
Xrepeater922 U$$2415/A1 VGND VGND VPWR VPWR U$$86/A1 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$729 final_adder.U$$712/A final_adder.U$$625/X final_adder.U$$609/X
+ VGND VGND VPWR VPWR final_adder.U$$729/X sky130_fd_sc_hd__a21o_2
XFILLER_99_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater933 input96/X VGND VGND VPWR VPWR U$$3646/A1 sky130_fd_sc_hd__buf_6
XFILLER_204_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater944 U$$4188/B1 VGND VGND VPWR VPWR U$$902/A1 sky130_fd_sc_hd__buf_6
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater955 U$$2955/A1 VGND VGND VPWR VPWR U$$3366/A1 sky130_fd_sc_hd__buf_4
Xrepeater966 input92/X VGND VGND VPWR VPWR U$$4460/A1 sky130_fd_sc_hd__buf_6
Xrepeater977 U$$2810/B1 VGND VGND VPWR VPWR U$$757/A1 sky130_fd_sc_hd__buf_6
XFILLER_204_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater988 U$$1209/B VGND VGND VPWR VPWR U$$1232/A sky130_fd_sc_hd__buf_12
Xrepeater999 input89/X VGND VGND VPWR VPWR U$$4178/B1 sky130_fd_sc_hd__buf_6
XFILLER_209_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3980 U$$3980/A U$$4012/B VGND VGND VPWR VPWR U$$3980/X sky130_fd_sc_hd__xor2_1
XU$$3991 U$$4402/A1 U$$4011/A2 U$$4402/B1 U$$4011/B2 VGND VGND VPWR VPWR U$$3992/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1915_1724 VGND VGND VPWR VPWR U$$1915_1724/HI U$$1915/B1 sky130_fd_sc_hd__conb_1
XFILLER_80_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_4_94_2 dadda_fa_4_94_2/A dadda_fa_4_94_2/B dadda_fa_4_94_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_95_0/CIN dadda_fa_5_94_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_118_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_87_1 dadda_fa_4_87_1/A dadda_fa_4_87_1/B dadda_fa_4_87_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/B dadda_fa_5_87_1/B sky130_fd_sc_hd__fa_1
XFILLER_134_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_64_0 dadda_fa_7_64_0/A dadda_fa_7_64_0/B dadda_fa_7_64_0/CIN VGND VGND
+ VPWR VPWR _361_/D _232_/D sky130_fd_sc_hd__fa_1
XFILLER_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput260 output260/A VGND VGND VPWR VPWR o[102] sky130_fd_sc_hd__buf_2
XFILLER_161_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput271 output271/A VGND VGND VPWR VPWR o[112] sky130_fd_sc_hd__buf_2
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput282 output282/A VGND VGND VPWR VPWR o[122] sky130_fd_sc_hd__buf_2
Xoutput293 output293/A VGND VGND VPWR VPWR o[17] sky130_fd_sc_hd__buf_2
XFILLER_47_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_1232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2008 U$$3102/B1 U$$2022/A2 U$$2967/B1 U$$2022/B2 VGND VGND VPWR VPWR U$$2009/A
+ sky130_fd_sc_hd__a22o_1
XU$$2019 U$$2019/A U$$2054/A VGND VGND VPWR VPWR U$$2019/X sky130_fd_sc_hd__xor2_1
XFILLER_55_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1307 U$$74/A1 U$$1311/A2 U$$1446/A1 U$$1307/B2 VGND VGND VPWR VPWR U$$1308/A sky130_fd_sc_hd__a22o_1
XFILLER_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1318 U$$1318/A U$$1366/B VGND VGND VPWR VPWR U$$1318/X sky130_fd_sc_hd__xor2_1
XFILLER_55_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1329 U$$96/A1 U$$1337/A2 U$$98/A1 U$$1337/B2 VGND VGND VPWR VPWR U$$1330/A sky130_fd_sc_hd__a22o_1
XFILLER_70_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_204_ _342_/CLK _204_/D VGND VGND VPWR VPWR _204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1101 final_adder.U$$178/B final_adder.U$$949/X VGND VGND VPWR VPWR
+ output359/A sky130_fd_sc_hd__xor2_1
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1112 final_adder.U$$166/A final_adder.U$$875/X VGND VGND VPWR VPWR
+ output371/A sky130_fd_sc_hd__xor2_1
XFILLER_184_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4107_1760 VGND VGND VPWR VPWR U$$4107_1760/HI U$$4107/B1 sky130_fd_sc_hd__conb_1
Xfinal_adder.U$$1123 final_adder.U$$156/B final_adder.U$$927/X VGND VGND VPWR VPWR
+ output383/A sky130_fd_sc_hd__xor2_1
XFILLER_183_243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1134 final_adder.U$$144/A final_adder.U$$853/X VGND VGND VPWR VPWR
+ output269/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1145 final_adder.U$$134/B final_adder.U$$905/X VGND VGND VPWR VPWR
+ output281/A sky130_fd_sc_hd__xor2_1
XFILLER_184_799 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_82_0 dadda_fa_3_82_0/A dadda_fa_3_82_0/B dadda_fa_3_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_0/B dadda_fa_4_82_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_180_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1018 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3210 U$$3210/A U$$3228/B VGND VGND VPWR VPWR U$$3210/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_111_0 U$$4485/X input142/X dadda_fa_4_111_0/CIN VGND VGND VPWR VPWR dadda_fa_5_112_0/A
+ dadda_fa_5_111_1/A sky130_fd_sc_hd__fa_1
XFILLER_24_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_44_5 dadda_fa_2_44_5/A dadda_fa_2_44_5/B dadda_fa_2_44_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_45_2/A dadda_fa_4_44_0/A sky130_fd_sc_hd__fa_1
XFILLER_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3221 U$$4178/B1 U$$3255/A2 U$$4045/A1 U$$3255/B2 VGND VGND VPWR VPWR U$$3222/A
+ sky130_fd_sc_hd__a22o_1
XU$$3232 U$$3232/A U$$3244/B VGND VGND VPWR VPWR U$$3232/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$14 _310_/Q _182_/Q VGND VGND VPWR VPWR final_adder.U$$241/A2 final_adder.U$$240/A
+ sky130_fd_sc_hd__ha_1
Xfinal_adder.U$$25 _321_/Q _193_/Q VGND VGND VPWR VPWR final_adder.U$$231/B1 final_adder.U$$230/B
+ sky130_fd_sc_hd__ha_1
XU$$3243 U$$3243/A1 U$$3155/X U$$3245/A1 U$$3156/X VGND VGND VPWR VPWR U$$3244/A sky130_fd_sc_hd__a22o_1
XFILLER_65_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3254 U$$3254/A U$$3256/B VGND VGND VPWR VPWR U$$3254/X sky130_fd_sc_hd__xor2_1
XFILLER_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3265 U$$251/A1 U$$3285/A2 U$$116/A1 U$$3285/B2 VGND VGND VPWR VPWR U$$3266/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$36 _332_/Q _204_/Q VGND VGND VPWR VPWR final_adder.U$$989/B1 final_adder.U$$218/A
+ sky130_fd_sc_hd__ha_1
XFILLER_19_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_37_4 U$$2342/X U$$2475/X input187/X VGND VGND VPWR VPWR dadda_fa_3_38_1/CIN
+ dadda_fa_3_37_3/CIN sky130_fd_sc_hd__fa_1
XU$$2520 U$$874/B1 U$$2542/A2 U$$741/A1 U$$2542/B2 VGND VGND VPWR VPWR U$$2521/A sky130_fd_sc_hd__a22o_1
XFILLER_111_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3276 U$$3276/A U$$3287/A VGND VGND VPWR VPWR U$$3276/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$47 _343_/Q _215_/Q VGND VGND VPWR VPWR final_adder.U$$209/B1 final_adder.U$$208/B
+ sky130_fd_sc_hd__ha_1
XU$$2531 U$$2531/A U$$2577/B VGND VGND VPWR VPWR U$$2531/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1084 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$58 _354_/Q _226_/Q VGND VGND VPWR VPWR final_adder.U$$967/B1 final_adder.U$$196/A
+ sky130_fd_sc_hd__ha_1
XU$$2542 U$$3499/B1 U$$2542/A2 U$$2955/A1 U$$2542/B2 VGND VGND VPWR VPWR U$$2543/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3287 U$$3287/A VGND VGND VPWR VPWR U$$3287/Y sky130_fd_sc_hd__inv_1
Xfinal_adder.U$$69 _365_/Q _237_/Q VGND VGND VPWR VPWR final_adder.U$$187/B1 final_adder.U$$186/B
+ sky130_fd_sc_hd__ha_1
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2553 U$$2553/A U$$2601/B VGND VGND VPWR VPWR U$$2553/X sky130_fd_sc_hd__xor2_1
XU$$3298 input76/X U$$3320/A2 U$$3300/A1 U$$3320/B2 VGND VGND VPWR VPWR U$$3299/A
+ sky130_fd_sc_hd__a22o_1
XU$$2564 U$$3112/A1 U$$2470/X U$$3114/A1 U$$2471/X VGND VGND VPWR VPWR U$$2565/A sky130_fd_sc_hd__a22o_1
XFILLER_181_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2575 U$$2575/A U$$2577/B VGND VGND VPWR VPWR U$$2575/X sky130_fd_sc_hd__xor2_1
XU$$1830 U$$1830/A U$$1832/B VGND VGND VPWR VPWR U$$1830/X sky130_fd_sc_hd__xor2_1
XU$$2586 U$$4365/B1 U$$2588/A2 U$$4095/A1 U$$2588/B2 VGND VGND VPWR VPWR U$$2587/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1841 U$$2113/B1 U$$1879/A2 U$$3348/B1 U$$1879/B2 VGND VGND VPWR VPWR U$$1842/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2597 U$$2597/A U$$2597/B VGND VGND VPWR VPWR U$$2597/X sky130_fd_sc_hd__xor2_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1852 U$$1852/A U$$1880/B VGND VGND VPWR VPWR U$$1852/X sky130_fd_sc_hd__xor2_1
XU$$1863 U$$2409/B1 U$$1869/A2 U$$3235/A1 U$$1869/B2 VGND VGND VPWR VPWR U$$1864/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1874 U$$1874/A U$$1878/B VGND VGND VPWR VPWR U$$1874/X sky130_fd_sc_hd__xor2_1
XU$$1885 U$$652/A1 U$$1915/A2 U$$517/A1 U$$1915/B2 VGND VGND VPWR VPWR U$$1886/A sky130_fd_sc_hd__a22o_1
XFILLER_159_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1896 U$$1896/A U$$1917/A VGND VGND VPWR VPWR U$$1896/X sky130_fd_sc_hd__xor2_1
XFILLER_159_251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_5_97_0 dadda_fa_5_97_0/A dadda_fa_5_97_0/B dadda_fa_5_97_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_98_0/A dadda_fa_6_97_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_174_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_803 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$515 final_adder.U$$514/B final_adder.U$$399/X final_adder.U$$391/X
+ VGND VGND VPWR VPWR final_adder.U$$515/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$526 final_adder.U$$534/B final_adder.U$$526/B VGND VGND VPWR VPWR
+ final_adder.U$$646/B sky130_fd_sc_hd__and2_1
Xrepeater730 U$$3517/B2 VGND VGND VPWR VPWR U$$3549/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$537 final_adder.U$$536/B final_adder.U$$421/X final_adder.U$$413/X
+ VGND VGND VPWR VPWR final_adder.U$$537/X sky130_fd_sc_hd__a21o_1
XTAP_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater741 U$$3293/X VGND VGND VPWR VPWR U$$3378/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$548 final_adder.U$$556/B final_adder.U$$548/B VGND VGND VPWR VPWR
+ final_adder.U$$668/B sky130_fd_sc_hd__and2_1
XTAP_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater752 U$$3019/X VGND VGND VPWR VPWR U$$3098/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$559 final_adder.U$$558/B final_adder.U$$443/X final_adder.U$$435/X
+ VGND VGND VPWR VPWR final_adder.U$$559/X sky130_fd_sc_hd__a21o_1
Xrepeater763 U$$2979/B2 VGND VGND VPWR VPWR U$$2967/B2 sky130_fd_sc_hd__buf_12
XU$$409 U$$409/A U$$410/A VGND VGND VPWR VPWR U$$409/X sky130_fd_sc_hd__xor2_1
Xrepeater774 U$$2796/B2 VGND VGND VPWR VPWR U$$2790/B2 sky130_fd_sc_hd__buf_4
Xrepeater785 U$$2691/B2 VGND VGND VPWR VPWR U$$2683/B2 sky130_fd_sc_hd__buf_6
XFILLER_84_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater796 U$$2558/B2 VGND VGND VPWR VPWR U$$2542/B2 sky130_fd_sc_hd__buf_8
XFILLER_72_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_916 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_811 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_938 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1309 U$$3377/B VGND VGND VPWR VPWR U$$3425/A sky130_fd_sc_hd__buf_6
XFILLER_101_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_106_1 U$$3943/X U$$4076/X U$$4209/X VGND VGND VPWR VPWR dadda_fa_4_107_0/CIN
+ dadda_fa_4_106_2/A sky130_fd_sc_hd__fa_1
XFILLER_69_23 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3011_1742 VGND VGND VPWR VPWR U$$3011_1742/HI U$$3011/B1 sky130_fd_sc_hd__conb_1
XFILLER_122_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_127_0 U$$4383/Y U$$4517/X input159/X VGND VGND VPWR VPWR dadda_fa_6_127_0/COUT
+ dadda_fa_7_127_0/CIN sky130_fd_sc_hd__fa_2
XFILLER_0_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_967 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_47_3 dadda_fa_3_47_3/A dadda_fa_3_47_3/B dadda_fa_3_47_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_48_1/B dadda_fa_4_47_2/CIN sky130_fd_sc_hd__fa_1
XU$$910 U$$910/A1 U$$918/A2 U$$912/A1 U$$918/B2 VGND VGND VPWR VPWR U$$911/A sky130_fd_sc_hd__a22o_1
XFILLER_29_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$921 U$$921/A U$$958/A VGND VGND VPWR VPWR U$$921/X sky130_fd_sc_hd__xor2_1
XFILLER_29_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$932 U$$932/A1 U$$938/A2 U$$932/B1 U$$938/B2 VGND VGND VPWR VPWR U$$933/A sky130_fd_sc_hd__a22o_1
XFILLER_91_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$943 U$$943/A U$$945/B VGND VGND VPWR VPWR U$$943/X sky130_fd_sc_hd__xor2_1
XFILLER_141_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$954 U$$954/A1 U$$826/X U$$956/A1 U$$827/X VGND VGND VPWR VPWR U$$955/A sky130_fd_sc_hd__a22o_1
XU$$965 U$$965/A1 U$$965/A2 U$$967/A1 U$$965/B2 VGND VGND VPWR VPWR U$$966/A sky130_fd_sc_hd__a22o_1
XU$$1104 U$$1515/A1 U$$1138/A2 U$$969/A1 U$$1138/B2 VGND VGND VPWR VPWR U$$1105/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_623 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$976 U$$976/A U$$980/B VGND VGND VPWR VPWR U$$976/X sky130_fd_sc_hd__xor2_1
XFILLER_16_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1115 U$$1115/A U$$1139/B VGND VGND VPWR VPWR U$$1115/X sky130_fd_sc_hd__xor2_1
XFILLER_203_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1126 U$$2357/B1 U$$1162/A2 U$$3594/A1 U$$1162/B2 VGND VGND VPWR VPWR U$$1127/A
+ sky130_fd_sc_hd__a22o_1
XU$$987 U$$987/A1 U$$999/A2 U$$987/B1 U$$999/B2 VGND VGND VPWR VPWR U$$988/A sky130_fd_sc_hd__a22o_1
XU$$1137 U$$1137/A U$$1137/B VGND VGND VPWR VPWR U$$1137/X sky130_fd_sc_hd__xor2_1
XU$$998 U$$998/A U$$998/B VGND VGND VPWR VPWR U$$998/X sky130_fd_sc_hd__xor2_1
XFILLER_188_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1148 U$$463/A1 U$$1162/A2 U$$54/A1 U$$1162/B2 VGND VGND VPWR VPWR U$$1149/A sky130_fd_sc_hd__a22o_1
XFILLER_188_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$1159 U$$1159/A U$$1195/B VGND VGND VPWR VPWR U$$1159/X sky130_fd_sc_hd__xor2_1
XFILLER_157_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_917 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1018 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_42_2 U$$2751/X U$$2884/X U$$2922/B VGND VGND VPWR VPWR dadda_fa_3_43_1/A
+ dadda_fa_3_42_3/A sky130_fd_sc_hd__fa_1
XFILLER_38_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3040 U$$3451/A1 U$$3124/A2 U$$28/A1 U$$3124/B2 VGND VGND VPWR VPWR U$$3041/A sky130_fd_sc_hd__a22o_1
Xclkbuf_3_4_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _239_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_208_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3051 U$$3051/A U$$3083/B VGND VGND VPWR VPWR U$$3051/X sky130_fd_sc_hd__xor2_1
XFILLER_187_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_35_1 U$$742/X U$$875/X U$$1008/X VGND VGND VPWR VPWR dadda_fa_3_36_0/CIN
+ dadda_fa_3_35_2/CIN sky130_fd_sc_hd__fa_1
XU$$3062 U$$3473/A1 U$$3098/A2 U$$4434/A1 U$$3098/B2 VGND VGND VPWR VPWR U$$3063/A
+ sky130_fd_sc_hd__a22o_1
XU$$3073 U$$3073/A U$$3077/B VGND VGND VPWR VPWR U$$3073/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_12_0 input160/X dadda_fa_5_12_0/B dadda_fa_5_12_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_6_13_0/A dadda_fa_6_12_0/CIN sky130_fd_sc_hd__fa_1
XU$$3084 U$$4454/A1 U$$3124/A2 U$$4456/A1 U$$3124/B2 VGND VGND VPWR VPWR U$$3085/A
+ sky130_fd_sc_hd__a22o_1
XU$$2350 U$$2350/A U$$2360/B VGND VGND VPWR VPWR U$$2350/X sky130_fd_sc_hd__xor2_1
XU$$3095 U$$3095/A U$$3151/A VGND VGND VPWR VPWR U$$3095/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_28_0 U$$63/X U$$196/X U$$329/X VGND VGND VPWR VPWR dadda_fa_3_29_1/CIN
+ dadda_fa_3_28_3/A sky130_fd_sc_hd__fa_1
XFILLER_34_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2361 U$$991/A1 U$$2417/A2 U$$2363/A1 U$$2417/B2 VGND VGND VPWR VPWR U$$2362/A
+ sky130_fd_sc_hd__a22o_1
XU$$2372 U$$2372/A U$$2380/B VGND VGND VPWR VPWR U$$2372/X sky130_fd_sc_hd__xor2_1
XFILLER_35_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2383 U$$3614/B1 U$$2417/A2 U$$3481/A1 U$$2417/B2 VGND VGND VPWR VPWR U$$2384/A
+ sky130_fd_sc_hd__a22o_1
XU$$2394 U$$2394/A U$$2442/B VGND VGND VPWR VPWR U$$2394/X sky130_fd_sc_hd__xor2_1
XU$$1660 U$$1932/B1 U$$1688/A2 U$$1799/A1 U$$1688/B2 VGND VGND VPWR VPWR U$$1661/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1671 U$$1671/A U$$1707/B VGND VGND VPWR VPWR U$$1671/X sky130_fd_sc_hd__xor2_1
XFILLER_195_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1682 U$$997/A1 U$$1688/A2 U$$997/B1 U$$1688/B2 VGND VGND VPWR VPWR U$$1683/A sky130_fd_sc_hd__a22o_1
XFILLER_61_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1693 U$$1693/A U$$1739/B VGND VGND VPWR VPWR U$$1693/X sky130_fd_sc_hd__xor2_1
XFILLER_148_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_87_4 U$$3240/X U$$3373/X U$$3506/X VGND VGND VPWR VPWR dadda_fa_2_88_4/B
+ dadda_fa_3_87_0/A sky130_fd_sc_hd__fa_1
XFILLER_39_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_170_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_57_2 dadda_fa_4_57_2/A dadda_fa_4_57_2/B dadda_fa_4_57_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_58_0/CIN dadda_fa_5_57_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_130_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$301 final_adder.U$$300/B final_adder.U$$175/X final_adder.U$$173/X
+ VGND VGND VPWR VPWR final_adder.U$$301/X sky130_fd_sc_hd__a21o_1
XTAP_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$312 final_adder.U$$314/B final_adder.U$$312/B VGND VGND VPWR VPWR
+ final_adder.U$$438/B sky130_fd_sc_hd__and2_1
XFILLER_170_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_945 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$323 final_adder.U$$322/B final_adder.U$$197/X final_adder.U$$195/X
+ VGND VGND VPWR VPWR final_adder.U$$323/X sky130_fd_sc_hd__a21o_1
XTAP_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$334 final_adder.U$$336/B final_adder.U$$334/B VGND VGND VPWR VPWR
+ final_adder.U$$460/B sky130_fd_sc_hd__and2_1
XTAP_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$345 final_adder.U$$344/B final_adder.U$$219/X final_adder.U$$217/X
+ VGND VGND VPWR VPWR final_adder.U$$345/X sky130_fd_sc_hd__a21o_1
XTAP_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$356 final_adder.U$$358/B final_adder.U$$356/B VGND VGND VPWR VPWR
+ final_adder.U$$482/B sky130_fd_sc_hd__and2_1
XTAP_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater560 U$$2252/A2 VGND VGND VPWR VPWR U$$2226/A2 sky130_fd_sc_hd__buf_6
Xdadda_fa_7_27_0 dadda_fa_7_27_0/A dadda_fa_7_27_0/B dadda_fa_7_27_0/CIN VGND VGND
+ VPWR VPWR _324_/D _195_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$367 final_adder.U$$366/B final_adder.U$$241/X final_adder.U$$239/X
+ VGND VGND VPWR VPWR final_adder.U$$367/X sky130_fd_sc_hd__a21o_1
XTAP_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$206 U$$206/A U$$212/B VGND VGND VPWR VPWR U$$206/X sky130_fd_sc_hd__xor2_1
Xrepeater571 U$$2169/A2 VGND VGND VPWR VPWR U$$2149/A2 sky130_fd_sc_hd__buf_6
XFILLER_85_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$378 final_adder.U$$378/A final_adder.U$$378/B VGND VGND VPWR VPWR
+ final_adder.U$$500/A sky130_fd_sc_hd__and2_1
XTAP_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater582 U$$1922/X VGND VGND VPWR VPWR U$$2040/A2 sky130_fd_sc_hd__buf_4
XU$$217 U$$80/A1 U$$217/A2 U$$82/A1 U$$217/B2 VGND VGND VPWR VPWR U$$218/A sky130_fd_sc_hd__a22o_1
XFILLER_73_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$389 final_adder.U$$388/B final_adder.U$$267/X final_adder.U$$263/X
+ VGND VGND VPWR VPWR final_adder.U$$389/X sky130_fd_sc_hd__a21o_1
XU$$228 U$$228/A U$$264/B VGND VGND VPWR VPWR U$$228/X sky130_fd_sc_hd__xor2_1
Xrepeater593 U$$1648/X VGND VGND VPWR VPWR U$$1736/A2 sky130_fd_sc_hd__buf_4
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$239 U$$787/A1 U$$243/A2 U$$926/A1 U$$243/B2 VGND VGND VPWR VPWR U$$240/A sky130_fd_sc_hd__a22o_1
XFILLER_72_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_1164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2609_1735 VGND VGND VPWR VPWR U$$2609_1735/HI U$$2609/A1 sky130_fd_sc_hd__conb_1
XFILLER_125_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1106 U$$3606/B1 VGND VGND VPWR VPWR U$$594/A1 sky130_fd_sc_hd__buf_4
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1080 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1117 input74/X VGND VGND VPWR VPWR U$$3878/B1 sky130_fd_sc_hd__buf_6
XFILLER_154_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1128 U$$4289/A1 VGND VGND VPWR VPWR U$$4426/A1 sky130_fd_sc_hd__buf_6
XFILLER_107_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1139 input71/X VGND VGND VPWR VPWR U$$312/A1 sky130_fd_sc_hd__buf_4
XFILLER_153_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_1170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_52_1 dadda_fa_3_52_1/A dadda_fa_3_52_1/B dadda_fa_3_52_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_0/CIN dadda_fa_4_52_2/A sky130_fd_sc_hd__fa_1
XFILLER_121_198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_68_1 U$$675/X U$$808/X U$$941/X VGND VGND VPWR VPWR dadda_fa_1_69_6/A
+ dadda_fa_1_68_7/CIN sky130_fd_sc_hd__fa_1
XFILLER_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_45_0 dadda_fa_3_45_0/A dadda_fa_3_45_0/B dadda_fa_3_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_0/B dadda_fa_4_45_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$740 U$$740/A U$$740/B VGND VGND VPWR VPWR U$$740/X sky130_fd_sc_hd__xor2_1
XFILLER_17_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$751 U$$888/A1 U$$759/A2 U$$890/A1 U$$759/B2 VGND VGND VPWR VPWR U$$752/A sky130_fd_sc_hd__a22o_1
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$762 U$$762/A U$$796/B VGND VGND VPWR VPWR U$$762/X sky130_fd_sc_hd__xor2_1
XU$$773 U$$910/A1 U$$783/A2 U$$773/B1 U$$783/B2 VGND VGND VPWR VPWR U$$774/A sky130_fd_sc_hd__a22o_1
XFILLER_205_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$784 U$$784/A U$$784/B VGND VGND VPWR VPWR U$$784/X sky130_fd_sc_hd__xor2_1
XFILLER_1_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$795 U$$930/B1 U$$805/A2 U$$932/B1 U$$805/B2 VGND VGND VPWR VPWR U$$796/A sky130_fd_sc_hd__a22o_1
XFILLER_91_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_ha_2_98_5 U$$4326/X U$$4459/X VGND VGND VPWR VPWR dadda_fa_3_99_2/B dadda_fa_4_98_0/A
+ sky130_fd_sc_hd__ha_1
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_185_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_7_102_0 dadda_fa_7_102_0/A dadda_fa_7_102_0/B dadda_fa_7_102_0/CIN VGND
+ VGND VPWR VPWR _399_/D _270_/D sky130_fd_sc_hd__fa_1
XFILLER_157_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_371 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_1 _327_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_97_3 U$$3526/X U$$3659/X U$$3792/X VGND VGND VPWR VPWR dadda_fa_3_98_1/B
+ dadda_fa_3_97_3/B sky130_fd_sc_hd__fa_1
Xrepeater1640 U$$2981/B1 VGND VGND VPWR VPWR U$$2709/A1 sky130_fd_sc_hd__buf_4
Xrepeater1651 U$$4488/A1 VGND VGND VPWR VPWR U$$789/A1 sky130_fd_sc_hd__buf_6
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1662 U$$783/B1 VGND VGND VPWR VPWR U$$920/B1 sky130_fd_sc_hd__buf_6
XFILLER_153_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1673 U$$4480/B1 VGND VGND VPWR VPWR U$$2016/A1 sky130_fd_sc_hd__buf_6
Xrepeater1684 input103/X VGND VGND VPWR VPWR U$$4478/B1 sky130_fd_sc_hd__buf_4
XFILLER_193_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1695 U$$3517/A1 VGND VGND VPWR VPWR U$$914/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_67_1 dadda_fa_5_67_1/A dadda_fa_5_67_1/B dadda_fa_5_67_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_68_0/B dadda_fa_7_67_0/A sky130_fd_sc_hd__fa_2
XFILLER_86_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_580 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_59_8 dadda_fa_1_59_8/A dadda_fa_1_59_8/B dadda_fa_1_59_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_60_3/A dadda_fa_3_59_0/A sky130_fd_sc_hd__fa_2
XFILLER_94_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_106_0 dadda_fa_2_106_0/A U$$3012/X U$$3145/X VGND VGND VPWR VPWR dadda_fa_3_107_3/B
+ dadda_fa_3_106_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_179_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2180 U$$2180/A input25/X VGND VGND VPWR VPWR U$$2180/X sky130_fd_sc_hd__xor2_1
XU$$2191 U$$2191/A VGND VGND VPWR VPWR U$$2191/Y sky130_fd_sc_hd__inv_1
XFILLER_210_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1490 U$$2449/A1 U$$1502/A2 U$$1764/B1 U$$1502/B2 VGND VGND VPWR VPWR U$$1491/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_1018 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_216 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_1_85_1 U$$1906/X U$$2039/X U$$2172/X VGND VGND VPWR VPWR dadda_fa_2_86_2/CIN
+ dadda_fa_2_85_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_116_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_62_0 dadda_fa_4_62_0/A dadda_fa_4_62_0/B dadda_fa_4_62_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/A dadda_fa_5_62_1/A sky130_fd_sc_hd__fa_1
XU$$6_1839 VGND VGND VPWR VPWR U$$6_1839/HI U$$6/A1 sky130_fd_sc_hd__conb_1
Xdadda_fa_1_78_0 U$$1227/X U$$1360/X U$$1493/X VGND VGND VPWR VPWR dadda_fa_2_79_0/B
+ dadda_fa_2_78_3/B sky130_fd_sc_hd__fa_1
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$120 _416_/Q _288_/Q VGND VGND VPWR VPWR final_adder.U$$905/B1 final_adder.U$$134/A
+ sky130_fd_sc_hd__ha_2
Xfinal_adder.U$$131 final_adder.U$$130/B final_adder.U$$901/B1 final_adder.U$$131/B1
+ VGND VGND VPWR VPWR final_adder.U$$131/X sky130_fd_sc_hd__a21o_1
XTAP_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3809 U$$3944/B1 U$$3813/A2 U$$3946/B1 U$$3813/B2 VGND VGND VPWR VPWR U$$3810/A
+ sky130_fd_sc_hd__a22o_1
XTAP_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$142 final_adder.U$$142/A final_adder.U$$142/B VGND VGND VPWR VPWR
+ final_adder.U$$270/B sky130_fd_sc_hd__and2_1
XTAP_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$153 final_adder.U$$152/B final_adder.U$$923/B1 final_adder.U$$153/B1
+ VGND VGND VPWR VPWR final_adder.U$$153/X sky130_fd_sc_hd__a21o_1
XTAP_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4388_1769 VGND VGND VPWR VPWR U$$4388_1769/HI U$$4388/A2 sky130_fd_sc_hd__conb_1
Xfinal_adder.U$$164 final_adder.U$$164/A final_adder.U$$164/B VGND VGND VPWR VPWR
+ final_adder.U$$292/B sky130_fd_sc_hd__and2_1
XTAP_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$175 final_adder.U$$174/B final_adder.U$$945/B1 final_adder.U$$175/B1
+ VGND VGND VPWR VPWR final_adder.U$$175/X sky130_fd_sc_hd__a21o_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1087 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$186 final_adder.U$$186/A final_adder.U$$186/B VGND VGND VPWR VPWR
+ final_adder.U$$314/B sky130_fd_sc_hd__and2_1
XTAP_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater390 U$$1083/A2 VGND VGND VPWR VPWR U$$1057/A2 sky130_fd_sc_hd__buf_4
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$197 final_adder.U$$196/B final_adder.U$$967/B1 final_adder.U$$197/B1
+ VGND VGND VPWR VPWR final_adder.U$$197/X sky130_fd_sc_hd__a21o_1
XTAP_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_452 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_383_ _385_/CLK _383_/D VGND VGND VPWR VPWR _383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1101 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_831 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_77_0 dadda_fa_6_77_0/A dadda_fa_6_77_0/B dadda_fa_6_77_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_78_0/B dadda_fa_7_77_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_147_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput160 c[12] VGND VGND VPWR VPWR input160/X sky130_fd_sc_hd__buf_4
XFILLER_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput171 c[22] VGND VGND VPWR VPWR input171/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$4447_1800 VGND VGND VPWR VPWR U$$4447_1800/HI U$$4447/B sky130_fd_sc_hd__conb_1
Xinput182 c[32] VGND VGND VPWR VPWR input182/X sky130_fd_sc_hd__buf_2
XFILLER_76_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput193 c[42] VGND VGND VPWR VPWR input193/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$570 U$$22/A1 U$$606/A2 U$$983/A1 U$$606/B2 VGND VGND VPWR VPWR U$$571/A sky130_fd_sc_hd__a22o_1
XU$$581 U$$581/A U$$607/B VGND VGND VPWR VPWR U$$581/X sky130_fd_sc_hd__xor2_1
XU$$592 U$$727/B1 U$$624/A2 U$$594/A1 U$$624/B2 VGND VGND VPWR VPWR U$$593/A sky130_fd_sc_hd__a22o_1
XFILLER_32_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_95_0 U$$2591/X U$$2724/X U$$2857/X VGND VGND VPWR VPWR dadda_fa_3_96_0/B
+ dadda_fa_3_95_2/B sky130_fd_sc_hd__fa_1
XFILLER_117_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1470 input127/X VGND VGND VPWR VPWR U$$3584/B1 sky130_fd_sc_hd__buf_8
XFILLER_99_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1481 U$$979/A1 VGND VGND VPWR VPWR U$$1799/B1 sky130_fd_sc_hd__buf_4
Xrepeater1492 U$$3283/B1 VGND VGND VPWR VPWR U$$3148/A1 sky130_fd_sc_hd__buf_4
XFILLER_87_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_71_7 dadda_fa_1_71_7/A dadda_fa_1_71_7/B dadda_fa_1_71_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_72_2/CIN dadda_fa_2_71_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_119_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_6 dadda_fa_1_64_6/A dadda_fa_1_64_6/B dadda_fa_1_64_6/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_2/B dadda_fa_2_64_5/B sky130_fd_sc_hd__fa_1
XFILLER_80_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_57_5 U$$3180/X U$$3313/X U$$3446/X VGND VGND VPWR VPWR dadda_fa_2_58_2/A
+ dadda_fa_2_57_5/A sky130_fd_sc_hd__fa_1
XFILLER_28_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_804 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1099 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_94_0 dadda_fa_7_94_0/A dadda_fa_7_94_0/B dadda_fa_7_94_0/CIN VGND VGND
+ VPWR VPWR _391_/D _262_/D sky130_fd_sc_hd__fa_2
XFILLER_183_639 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_920 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4307 U$$4307/A1 U$$4381/A2 U$$4309/A1 U$$4381/B2 VGND VGND VPWR VPWR U$$4308/A
+ sky130_fd_sc_hd__a22o_1
XU$$4318 U$$4318/A U$$4330/B VGND VGND VPWR VPWR U$$4318/X sky130_fd_sc_hd__xor2_1
XFILLER_19_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4329 U$$4466/A1 U$$4349/A2 U$$4466/B1 U$$4349/B2 VGND VGND VPWR VPWR U$$4330/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3606 U$$3878/B1 U$$3606/A2 U$$3606/B1 U$$3606/B2 VGND VGND VPWR VPWR U$$3607/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3617 U$$3617/A U$$3623/B VGND VGND VPWR VPWR U$$3617/X sky130_fd_sc_hd__xor2_1
XFILLER_19_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3628 U$$4311/B1 U$$3566/X U$$4176/B1 U$$3567/X VGND VGND VPWR VPWR U$$3629/A sky130_fd_sc_hd__a22o_1
XU$$3639 U$$3639/A U$$3643/B VGND VGND VPWR VPWR U$$3639/X sky130_fd_sc_hd__xor2_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2905 U$$28/A1 U$$2919/A2 U$$30/A1 U$$2919/B2 VGND VGND VPWR VPWR U$$2906/A sky130_fd_sc_hd__a22o_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2916 U$$2916/A U$$2920/B VGND VGND VPWR VPWR U$$2916/X sky130_fd_sc_hd__xor2_1
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2927 U$$461/A1 U$$2949/A2 U$$4297/B1 U$$2949/B2 VGND VGND VPWR VPWR U$$2928/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 _200_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2938 U$$2938/A U$$2968/B VGND VGND VPWR VPWR U$$2938/X sky130_fd_sc_hd__xor2_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2949 U$$2949/A1 U$$2949/A2 U$$2951/A1 U$$2949/B2 VGND VGND VPWR VPWR U$$2950/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_3_22_2 U$$1115/X U$$1248/X U$$1381/X VGND VGND VPWR VPWR dadda_fa_4_23_1/A
+ dadda_fa_4_22_2/B sky130_fd_sc_hd__fa_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_243 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 input109/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 U$$1877/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_366_ _367_/CLK _366_/D VGND VGND VPWR VPWR _366_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4477_1815 VGND VGND VPWR VPWR U$$4477_1815/HI U$$4477/B sky130_fd_sc_hd__conb_1
XFILLER_158_168 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_297_ _304_/CLK _297_/D VGND VGND VPWR VPWR _297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_74_5 dadda_fa_2_74_5/A dadda_fa_2_74_5/B dadda_fa_2_74_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_75_2/A dadda_fa_4_74_0/A sky130_fd_sc_hd__fa_1
XFILLER_111_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_67_4 dadda_fa_2_67_4/A dadda_fa_2_67_4/B dadda_fa_2_67_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_1/CIN dadda_fa_3_67_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_110_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_989 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_973 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_945 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_5_104_1 dadda_fa_5_104_1/A dadda_fa_5_104_1/B dadda_fa_5_104_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_105_0/B dadda_fa_7_104_0/A sky130_fd_sc_hd__fa_2
XFILLER_145_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_472 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_62_3 U$$3589/X U$$3722/X U$$3855/X VGND VGND VPWR VPWR dadda_fa_2_63_1/B
+ dadda_fa_2_62_4/B sky130_fd_sc_hd__fa_1
XFILLER_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_55_2 U$$1580/X U$$1713/X U$$1846/X VGND VGND VPWR VPWR dadda_fa_2_56_1/A
+ dadda_fa_2_55_4/A sky130_fd_sc_hd__fa_1
XFILLER_170_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_32_1 dadda_fa_4_32_1/A dadda_fa_4_32_1/B dadda_fa_4_32_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/B dadda_fa_5_32_1/B sky130_fd_sc_hd__fa_1
XFILLER_103_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_48_1 U$$502/X U$$635/X U$$768/X VGND VGND VPWR VPWR dadda_fa_2_49_1/B
+ dadda_fa_2_48_4/A sky130_fd_sc_hd__fa_1
XFILLER_103_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_25_0 dadda_fa_4_25_0/A dadda_fa_4_25_0/B dadda_fa_4_25_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/A dadda_fa_5_25_1/A sky130_fd_sc_hd__fa_1
XFILLER_167_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_220_ _351_/CLK _220_/D VGND VGND VPWR VPWR _220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_948 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_174_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_77_3 dadda_fa_3_77_3/A dadda_fa_3_77_3/B dadda_fa_3_77_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_78_1/B dadda_fa_4_77_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4104 U$$4104/A input55/X VGND VGND VPWR VPWR U$$4104/X sky130_fd_sc_hd__xor2_1
XFILLER_24_1230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4115 U$$4113/B input55/X input57/X U$$4110/Y VGND VGND VPWR VPWR U$$4115/X sky130_fd_sc_hd__a22o_2
XFILLER_78_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4126 U$$4400/A1 U$$4144/A2 U$$4402/A1 U$$4144/B2 VGND VGND VPWR VPWR U$$4127/A
+ sky130_fd_sc_hd__a22o_1
XU$$4137 U$$4137/A U$$4165/B VGND VGND VPWR VPWR U$$4137/X sky130_fd_sc_hd__xor2_1
XU$$3403 U$$3403/A U$$3424/A VGND VGND VPWR VPWR U$$3403/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_14_0 U$$35/X U$$168/X VGND VGND VPWR VPWR dadda_fa_4_15_2/B dadda_ha_3_14_0/SUM
+ sky130_fd_sc_hd__ha_1
XU$$4148 input71/X U$$4188/A2 input72/X U$$4188/B2 VGND VGND VPWR VPWR U$$4149/A sky130_fd_sc_hd__a22o_1
XU$$3414 U$$3414/A1 U$$3416/A2 U$$3414/B1 U$$3416/B2 VGND VGND VPWR VPWR U$$3415/A
+ sky130_fd_sc_hd__a22o_1
XU$$4159 U$$4159/A U$$4165/B VGND VGND VPWR VPWR U$$4159/X sky130_fd_sc_hd__xor2_1
XU$$3425 U$$3425/A VGND VGND VPWR VPWR U$$3425/Y sky130_fd_sc_hd__inv_1
XFILLER_92_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3436 U$$3436/A U$$3528/B VGND VGND VPWR VPWR U$$3436/X sky130_fd_sc_hd__xor2_1
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2702 U$$2702/A U$$2710/B VGND VGND VPWR VPWR U$$2702/X sky130_fd_sc_hd__xor2_1
XFILLER_80_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3447 U$$3447/A1 U$$3453/A2 U$$3584/B1 U$$3453/B2 VGND VGND VPWR VPWR U$$3448/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3458 U$$3458/A U$$3480/B VGND VGND VPWR VPWR U$$3458/X sky130_fd_sc_hd__xor2_1
XU$$2713 U$$4494/A1 U$$2737/A2 U$$2715/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2714/A
+ sky130_fd_sc_hd__a22o_1
XU$$2724 U$$2724/A U$$2736/B VGND VGND VPWR VPWR U$$2724/X sky130_fd_sc_hd__xor2_1
XU$$3469 U$$4428/A1 U$$3503/A2 U$$4430/A1 U$$3503/B2 VGND VGND VPWR VPWR U$$3470/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2735 U$$3281/B1 U$$2735/A2 U$$3148/A1 U$$2735/B2 VGND VGND VPWR VPWR U$$2736/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2746 U$$2746/A1 U$$2796/A2 U$$3159/A1 U$$2796/B2 VGND VGND VPWR VPWR U$$2747/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2757 U$$2757/A U$$2797/B VGND VGND VPWR VPWR U$$2757/X sky130_fd_sc_hd__xor2_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2768 U$$711/B1 U$$2782/A2 U$$578/A1 U$$2782/B2 VGND VGND VPWR VPWR U$$2769/A sky130_fd_sc_hd__a22o_1
XU$$2779 U$$2779/A U$$2783/B VGND VGND VPWR VPWR U$$2779/X sky130_fd_sc_hd__xor2_1
XFILLER_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1001 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_418_ _419_/CLK _418_/D VGND VGND VPWR VPWR _418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_349_ _351_/CLK _349_/D VGND VGND VPWR VPWR _349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_72_2 dadda_fa_2_72_2/A dadda_fa_2_72_2/B dadda_fa_2_72_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/A dadda_fa_3_72_3/A sky130_fd_sc_hd__fa_1
XFILLER_130_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_65_1 dadda_fa_2_65_1/A dadda_fa_2_65_1/B dadda_fa_2_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_0/CIN dadda_fa_3_65_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_9_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_818 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater901 U$$4512/B2 VGND VGND VPWR VPWR U$$4498/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$708 final_adder.U$$708/A final_adder.U$$708/B VGND VGND VPWR VPWR
+ final_adder.U$$788/A sky130_fd_sc_hd__and2_1
Xrepeater912 U$$2069/A1 VGND VGND VPWR VPWR U$$836/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_96_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$719 final_adder.U$$718/B final_adder.U$$615/X final_adder.U$$599/X
+ VGND VGND VPWR VPWR final_adder.U$$719/X sky130_fd_sc_hd__a21o_1
Xdadda_fa_5_42_0 dadda_fa_5_42_0/A dadda_fa_5_42_0/B dadda_fa_5_42_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_43_0/A dadda_fa_6_42_0/CIN sky130_fd_sc_hd__fa_1
Xrepeater923 U$$3235/B1 VGND VGND VPWR VPWR U$$2415/A1 sky130_fd_sc_hd__buf_12
Xrepeater934 input96/X VGND VGND VPWR VPWR U$$4466/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_58_0 dadda_fa_2_58_0/A dadda_fa_2_58_0/B dadda_fa_2_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_0/B dadda_fa_3_58_2/B sky130_fd_sc_hd__fa_1
Xrepeater945 U$$3366/B1 VGND VGND VPWR VPWR U$$763/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_83_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater956 input93/X VGND VGND VPWR VPWR U$$2955/A1 sky130_fd_sc_hd__buf_8
Xrepeater967 U$$2951/A1 VGND VGND VPWR VPWR U$$74/A1 sky130_fd_sc_hd__buf_4
XFILLER_209_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater978 U$$2810/B1 VGND VGND VPWR VPWR U$$894/A1 sky130_fd_sc_hd__buf_6
Xrepeater989 U$$1205/B VGND VGND VPWR VPWR U$$1195/B sky130_fd_sc_hd__buf_6
XFILLER_204_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_873 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3970 U$$4242/B1 U$$3970/A2 U$$3970/B1 U$$3970/B2 VGND VGND VPWR VPWR U$$3971/A
+ sky130_fd_sc_hd__a22o_1
XU$$3981 U$$4392/A1 U$$4011/A2 U$$4394/A1 U$$4011/B2 VGND VGND VPWR VPWR U$$3982/A
+ sky130_fd_sc_hd__a22o_1
XU$$3992 U$$3992/A U$$4012/B VGND VGND VPWR VPWR U$$3992/X sky130_fd_sc_hd__xor2_1
XFILLER_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1025 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_1167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_948 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_87_2 dadda_fa_4_87_2/A dadda_fa_4_87_2/B dadda_fa_4_87_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_88_0/CIN dadda_fa_5_87_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput261 output261/A VGND VGND VPWR VPWR o[103] sky130_fd_sc_hd__buf_2
Xdadda_fa_7_57_0 dadda_fa_7_57_0/A dadda_fa_7_57_0/B dadda_fa_7_57_0/CIN VGND VGND
+ VPWR VPWR _354_/D _225_/D sky130_fd_sc_hd__fa_1
Xoutput272 output272/A VGND VGND VPWR VPWR o[113] sky130_fd_sc_hd__buf_2
XFILLER_161_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput283 output283/A VGND VGND VPWR VPWR o[123] sky130_fd_sc_hd__buf_2
XFILLER_82_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput294 output294/A VGND VGND VPWR VPWR o[18] sky130_fd_sc_hd__buf_2
XFILLER_173_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_60_0 U$$1989/X U$$2122/X U$$2255/X VGND VGND VPWR VPWR dadda_fa_2_61_0/B
+ dadda_fa_2_60_3/B sky130_fd_sc_hd__fa_1
XFILLER_75_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2009 U$$2009/A U$$2009/B VGND VGND VPWR VPWR U$$2009/X sky130_fd_sc_hd__xor2_1
XFILLER_62_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1308 U$$1308/A U$$1316/B VGND VGND VPWR VPWR U$$1308/X sky130_fd_sc_hd__xor2_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1319 U$$3922/A1 U$$1353/A2 U$$3922/B1 U$$1355/B2 VGND VGND VPWR VPWR U$$1320/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_943 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_203_ _337_/CLK _203_/D VGND VGND VPWR VPWR _203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_965 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_639 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1102 final_adder.U$$176/A final_adder.U$$885/X VGND VGND VPWR VPWR
+ output360/A sky130_fd_sc_hd__xor2_1
XFILLER_12_998 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1113 final_adder.U$$166/B final_adder.U$$937/X VGND VGND VPWR VPWR
+ output372/A sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$1124 final_adder.U$$154/A final_adder.U$$863/X VGND VGND VPWR VPWR
+ output258/A sky130_fd_sc_hd__xor2_2
XFILLER_172_907 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1135 final_adder.U$$144/B final_adder.U$$915/X VGND VGND VPWR VPWR
+ output270/A sky130_fd_sc_hd__xor2_1
XFILLER_183_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1146 final_adder.U$$132/A final_adder.U$$841/X VGND VGND VPWR VPWR
+ output282/A sky130_fd_sc_hd__xor2_1
XFILLER_171_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_1171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_82_1 dadda_fa_3_82_1/A dadda_fa_3_82_1/B dadda_fa_3_82_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_0/CIN dadda_fa_4_82_2/A sky130_fd_sc_hd__fa_1
XFILLER_48_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_75_0 dadda_fa_3_75_0/A dadda_fa_3_75_0/B dadda_fa_3_75_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_0/B dadda_fa_4_75_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3200 U$$3200/A U$$3242/B VGND VGND VPWR VPWR U$$3200/X sky130_fd_sc_hd__xor2_1
XFILLER_65_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3211 U$$3485/A1 U$$3229/A2 U$$3211/B1 U$$3227/B2 VGND VGND VPWR VPWR U$$3212/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_111_1 dadda_fa_4_111_1/A dadda_fa_4_111_1/B dadda_fa_4_111_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_112_0/B dadda_fa_5_111_1/B sky130_fd_sc_hd__fa_1
XFILLER_93_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3222 U$$3222/A U$$3256/B VGND VGND VPWR VPWR U$$3222/X sky130_fd_sc_hd__xor2_1
XFILLER_24_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3233 U$$3368/B1 U$$3241/A2 U$$3235/A1 U$$3241/B2 VGND VGND VPWR VPWR U$$3234/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$15 _311_/Q _183_/Q VGND VGND VPWR VPWR final_adder.U$$241/B1 final_adder.U$$240/B
+ sky130_fd_sc_hd__ha_1
XFILLER_0_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3244 U$$3244/A U$$3244/B VGND VGND VPWR VPWR U$$3244/X sky130_fd_sc_hd__xor2_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$26 _322_/Q _194_/Q VGND VGND VPWR VPWR final_adder.U$$999/B1 final_adder.U$$228/A
+ sky130_fd_sc_hd__ha_1
XU$$3255 U$$3801/B1 U$$3255/A2 U$$517/A1 U$$3255/B2 VGND VGND VPWR VPWR U$$3256/A
+ sky130_fd_sc_hd__a22o_1
XU$$2510 U$$4015/B1 U$$2596/A2 U$$3880/B1 U$$2596/B2 VGND VGND VPWR VPWR U$$2511/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_104_0 dadda_fa_4_104_0/A dadda_fa_4_104_0/B dadda_fa_4_104_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/A dadda_fa_5_104_1/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$37 _333_/Q _205_/Q VGND VGND VPWR VPWR final_adder.U$$219/B1 final_adder.U$$218/B
+ sky130_fd_sc_hd__ha_1
Xdadda_fa_2_37_5 dadda_fa_2_37_5/A dadda_fa_2_37_5/B dadda_fa_2_37_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_38_2/A dadda_fa_4_37_0/A sky130_fd_sc_hd__fa_1
XU$$3266 U$$3266/A U$$3286/B VGND VGND VPWR VPWR U$$3266/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$48 _344_/Q _216_/Q VGND VGND VPWR VPWR final_adder.U$$977/B1 final_adder.U$$206/A
+ sky130_fd_sc_hd__ha_1
XFILLER_19_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2521 U$$2521/A U$$2543/B VGND VGND VPWR VPWR U$$2521/X sky130_fd_sc_hd__xor2_1
XFILLER_206_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3277 U$$3551/A1 U$$3277/A2 input121/X U$$3277/B2 VGND VGND VPWR VPWR U$$3278/A
+ sky130_fd_sc_hd__a22o_1
XU$$2532 U$$4176/A1 U$$2576/A2 U$$3902/B1 U$$2576/B2 VGND VGND VPWR VPWR U$$2533/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$59 _355_/Q _227_/Q VGND VGND VPWR VPWR final_adder.U$$197/B1 final_adder.U$$196/B
+ sky130_fd_sc_hd__ha_1
XU$$2543 U$$2543/A U$$2543/B VGND VGND VPWR VPWR U$$2543/X sky130_fd_sc_hd__xor2_1
XU$$3288 U$$3288/A VGND VGND VPWR VPWR U$$3288/Y sky130_fd_sc_hd__inv_1
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2554 U$$3922/B1 U$$2588/A2 U$$3787/B1 U$$2588/B2 VGND VGND VPWR VPWR U$$2555/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3299 U$$3299/A U$$3321/B VGND VGND VPWR VPWR U$$3299/X sky130_fd_sc_hd__xor2_1
XFILLER_181_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1820 U$$1820/A U$$1820/B VGND VGND VPWR VPWR U$$1820/X sky130_fd_sc_hd__xor2_1
XFILLER_55_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2565 U$$2565/A U$$2603/A VGND VGND VPWR VPWR U$$2565/X sky130_fd_sc_hd__xor2_1
XFILLER_185_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1831 U$$2925/B1 U$$1831/A2 U$$3612/B1 U$$1831/B2 VGND VGND VPWR VPWR U$$1832/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2576 U$$2711/B1 U$$2576/A2 U$$934/A1 U$$2576/B2 VGND VGND VPWR VPWR U$$2577/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2587 U$$2587/A U$$2602/A VGND VGND VPWR VPWR U$$2587/X sky130_fd_sc_hd__xor2_1
XU$$1842 U$$1842/A U$$1880/B VGND VGND VPWR VPWR U$$1842/X sky130_fd_sc_hd__xor2_1
XU$$2598 U$$3281/B1 U$$2600/A2 U$$3148/A1 U$$2600/B2 VGND VGND VPWR VPWR U$$2599/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1853 U$$2949/A1 U$$1879/A2 U$$483/B1 U$$1879/B2 VGND VGND VPWR VPWR U$$1854/A
+ sky130_fd_sc_hd__a22o_1
XU$$1864 U$$1864/A U$$1870/B VGND VGND VPWR VPWR U$$1864/X sky130_fd_sc_hd__xor2_1
XU$$1875 U$$2834/A1 U$$1877/A2 U$$2425/A1 U$$1877/B2 VGND VGND VPWR VPWR U$$1876/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1886 U$$1886/A U$$1917/A VGND VGND VPWR VPWR U$$1886/X sky130_fd_sc_hd__xor2_1
XFILLER_61_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1897 U$$2582/A1 U$$1915/A2 U$$4502/A1 U$$1915/B2 VGND VGND VPWR VPWR U$$1898/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_97_1 dadda_fa_5_97_1/A dadda_fa_5_97_1/B dadda_fa_5_97_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_98_0/B dadda_fa_7_97_0/A sky130_fd_sc_hd__fa_1
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$505 final_adder.U$$500/A final_adder.U$$255/X final_adder.U$$379/X
+ VGND VGND VPWR VPWR final_adder.U$$505/X sky130_fd_sc_hd__a21o_2
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$516 final_adder.U$$524/B final_adder.U$$516/B VGND VGND VPWR VPWR
+ final_adder.U$$636/B sky130_fd_sc_hd__and2_1
Xrepeater720 U$$3644/B2 VGND VGND VPWR VPWR U$$3660/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$527 final_adder.U$$526/B final_adder.U$$411/X final_adder.U$$403/X
+ VGND VGND VPWR VPWR final_adder.U$$527/X sky130_fd_sc_hd__a21o_1
Xrepeater731 U$$3517/B2 VGND VGND VPWR VPWR U$$3559/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$538 final_adder.U$$546/B final_adder.U$$538/B VGND VGND VPWR VPWR
+ final_adder.U$$658/B sky130_fd_sc_hd__and2_1
XTAP_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater742 U$$3227/B2 VGND VGND VPWR VPWR U$$3187/B2 sky130_fd_sc_hd__buf_4
Xfinal_adder.U$$549 final_adder.U$$548/B final_adder.U$$433/X final_adder.U$$425/X
+ VGND VGND VPWR VPWR final_adder.U$$549/X sky130_fd_sc_hd__a21o_1
Xrepeater753 U$$3132/B2 VGND VGND VPWR VPWR U$$3124/B2 sky130_fd_sc_hd__buf_6
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater764 U$$2882/X VGND VGND VPWR VPWR U$$2979/B2 sky130_fd_sc_hd__buf_4
XFILLER_84_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater775 U$$2810/B2 VGND VGND VPWR VPWR U$$2796/B2 sky130_fd_sc_hd__buf_4
XFILLER_44_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater786 U$$2711/B2 VGND VGND VPWR VPWR U$$2691/B2 sky130_fd_sc_hd__buf_6
XFILLER_77_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater797 U$$2471/X VGND VGND VPWR VPWR U$$2558/B2 sky130_fd_sc_hd__buf_6
XFILLER_71_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4490 U$$4490/A1 U$$4388/X U$$4492/A1 U$$4494/B2 VGND VGND VPWR VPWR U$$4491/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_915 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_92_0 dadda_fa_4_92_0/A dadda_fa_4_92_0/B dadda_fa_4_92_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/A dadda_fa_5_92_1/A sky130_fd_sc_hd__fa_1
XFILLER_158_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_106_2 U$$4342/X U$$4475/X input136/X VGND VGND VPWR VPWR dadda_fa_4_107_1/A
+ dadda_fa_4_106_2/B sky130_fd_sc_hd__fa_1
XFILLER_134_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_675 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_919 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$900 U$$78/A1 U$$906/A2 U$$80/A1 U$$906/B2 VGND VGND VPWR VPWR U$$901/A sky130_fd_sc_hd__a22o_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$911 U$$911/A U$$919/B VGND VGND VPWR VPWR U$$911/X sky130_fd_sc_hd__xor2_1
XFILLER_28_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$922 U$$98/B1 U$$950/A2 U$$924/A1 U$$950/B2 VGND VGND VPWR VPWR U$$923/A sky130_fd_sc_hd__a22o_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$933 U$$933/A U$$945/B VGND VGND VPWR VPWR U$$933/X sky130_fd_sc_hd__xor2_1
XFILLER_44_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$944 U$$944/A1 U$$950/A2 U$$944/B1 U$$950/B2 VGND VGND VPWR VPWR U$$945/A sky130_fd_sc_hd__a22o_1
XU$$955 U$$955/A U$$958/A VGND VGND VPWR VPWR U$$955/X sky130_fd_sc_hd__xor2_1
XU$$1105 U$$1105/A U$$1139/B VGND VGND VPWR VPWR U$$1105/X sky130_fd_sc_hd__xor2_1
XU$$966 U$$966/A U$$968/B VGND VGND VPWR VPWR U$$966/X sky130_fd_sc_hd__xor2_1
XFILLER_204_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1116 U$$1799/B1 U$$1136/A2 U$$981/A1 U$$1136/B2 VGND VGND VPWR VPWR U$$1117/A
+ sky130_fd_sc_hd__a22o_1
XU$$977 U$$18/A1 U$$979/A2 U$$979/A1 U$$979/B2 VGND VGND VPWR VPWR U$$978/A sky130_fd_sc_hd__a22o_1
XU$$1127 U$$1127/A U$$1195/B VGND VGND VPWR VPWR U$$1127/X sky130_fd_sc_hd__xor2_1
XU$$988 U$$988/A U$$996/B VGND VGND VPWR VPWR U$$988/X sky130_fd_sc_hd__xor2_1
XU$$999 U$$999/A1 U$$999/A2 U$$42/A1 U$$999/B2 VGND VGND VPWR VPWR U$$999/X sky130_fd_sc_hd__a22o_1
XU$$1138 U$$179/A1 U$$1138/A2 U$$866/A1 U$$1138/B2 VGND VGND VPWR VPWR U$$1139/A sky130_fd_sc_hd__a22o_1
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1149 U$$1149/A U$$1187/B VGND VGND VPWR VPWR U$$1149/X sky130_fd_sc_hd__xor2_1
XFILLER_43_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_870 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_929 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_642 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_984 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_2_29_3 U$$1262/X U$$1395/X VGND VGND VPWR VPWR dadda_fa_3_30_2/B dadda_fa_4_29_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_1147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_42_3 input193/X dadda_fa_2_42_3/B dadda_fa_2_42_3/CIN VGND VGND VPWR VPWR
+ dadda_fa_3_43_1/B dadda_fa_3_42_3/B sky130_fd_sc_hd__fa_1
XFILLER_54_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1248 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3030 input109/X U$$3082/A2 U$$3578/B1 U$$3082/B2 VGND VGND VPWR VPWR U$$3031/A
+ sky130_fd_sc_hd__a22o_1
XU$$3041 U$$3041/A U$$3125/B VGND VGND VPWR VPWR U$$3041/X sky130_fd_sc_hd__xor2_1
XFILLER_82_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3052 U$$4011/A1 U$$3082/A2 U$$4011/B1 U$$3082/B2 VGND VGND VPWR VPWR U$$3053/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3063 U$$3063/A U$$3077/B VGND VGND VPWR VPWR U$$3063/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_2 U$$1141/X U$$1274/X U$$1407/X VGND VGND VPWR VPWR dadda_fa_3_36_1/A
+ dadda_fa_3_35_3/A sky130_fd_sc_hd__fa_1
XU$$3074 U$$3485/A1 U$$3098/A2 U$$610/A1 U$$3098/B2 VGND VGND VPWR VPWR U$$3075/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2340 U$$2340/A U$$2366/B VGND VGND VPWR VPWR U$$2340/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_5_12_1 dadda_fa_5_12_1/A dadda_fa_5_12_1/B dadda_ha_4_12_2/SUM VGND VGND
+ VPWR VPWR dadda_fa_6_13_0/B dadda_fa_7_12_0/A sky130_fd_sc_hd__fa_1
XU$$3085 U$$3085/A U$$3125/B VGND VGND VPWR VPWR U$$3085/X sky130_fd_sc_hd__xor2_1
XFILLER_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2351 U$$2625/A1 U$$2359/A2 U$$2625/B1 U$$2359/B2 VGND VGND VPWR VPWR U$$2352/A
+ sky130_fd_sc_hd__a22o_1
Xdadda_fa_2_28_1 U$$462/X U$$595/X U$$728/X VGND VGND VPWR VPWR dadda_fa_3_29_2/A
+ dadda_fa_3_28_3/B sky130_fd_sc_hd__fa_1
XU$$3096 U$$3644/A1 U$$3018/X U$$3644/B1 U$$3019/X VGND VGND VPWR VPWR U$$3097/A sky130_fd_sc_hd__a22o_1
XFILLER_50_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2362 U$$2362/A U$$2366/B VGND VGND VPWR VPWR U$$2362/X sky130_fd_sc_hd__xor2_1
XU$$2373 U$$4015/B1 U$$2463/A2 U$$3880/B1 U$$2463/B2 VGND VGND VPWR VPWR U$$2374/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2384 U$$2384/A U$$2426/B VGND VGND VPWR VPWR U$$2384/X sky130_fd_sc_hd__xor2_1
XFILLER_62_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1650 U$$1650/A1 U$$1696/A2 U$$2198/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1651/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2395 U$$3078/B1 U$$2403/A2 U$$890/A1 U$$2403/B2 VGND VGND VPWR VPWR U$$2396/A
+ sky130_fd_sc_hd__a22o_1
XU$$1661 U$$1661/A U$$1689/B VGND VGND VPWR VPWR U$$1661/X sky130_fd_sc_hd__xor2_1
XU$$1672 U$$850/A1 U$$1706/A2 U$$850/B1 U$$1706/B2 VGND VGND VPWR VPWR U$$1673/A sky130_fd_sc_hd__a22o_1
XFILLER_148_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1683 U$$1683/A U$$1689/B VGND VGND VPWR VPWR U$$1683/X sky130_fd_sc_hd__xor2_1
XU$$1694 U$$598/A1 U$$1746/A2 U$$463/A1 U$$1746/B2 VGND VGND VPWR VPWR U$$1695/A sky130_fd_sc_hd__a22o_1
XFILLER_148_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$302 final_adder.U$$304/B final_adder.U$$302/B VGND VGND VPWR VPWR
+ final_adder.U$$428/B sky130_fd_sc_hd__and2_1
XTAP_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$313 final_adder.U$$312/B final_adder.U$$187/X final_adder.U$$185/X
+ VGND VGND VPWR VPWR final_adder.U$$313/X sky130_fd_sc_hd__a21o_1
XTAP_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$324 final_adder.U$$326/B final_adder.U$$324/B VGND VGND VPWR VPWR
+ final_adder.U$$450/B sky130_fd_sc_hd__and2_1
XFILLER_58_957 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$335 final_adder.U$$334/B final_adder.U$$209/X final_adder.U$$207/X
+ VGND VGND VPWR VPWR final_adder.U$$335/X sky130_fd_sc_hd__a21o_1
XTAP_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$346 final_adder.U$$348/B final_adder.U$$346/B VGND VGND VPWR VPWR
+ final_adder.U$$472/B sky130_fd_sc_hd__and2_1
XTAP_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater550 U$$2470/X VGND VGND VPWR VPWR U$$2558/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$357 final_adder.U$$356/B final_adder.U$$231/X final_adder.U$$229/X
+ VGND VGND VPWR VPWR final_adder.U$$357/X sky130_fd_sc_hd__a21o_1
XTAP_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater561 U$$2302/A2 VGND VGND VPWR VPWR U$$2252/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_84_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$368 final_adder.U$$370/B final_adder.U$$368/B VGND VGND VPWR VPWR
+ final_adder.U$$494/B sky130_fd_sc_hd__and2_1
XTAP_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$207 U$$70/A1 U$$259/A2 U$$72/A1 U$$259/B2 VGND VGND VPWR VPWR U$$208/A sky130_fd_sc_hd__a22o_1
Xrepeater572 U$$2183/A2 VGND VGND VPWR VPWR U$$2189/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$379 final_adder.U$$378/B final_adder.U$$253/X final_adder.U$$251/X
+ VGND VGND VPWR VPWR final_adder.U$$379/X sky130_fd_sc_hd__a21o_1
XU$$218 U$$218/A U$$218/B VGND VGND VPWR VPWR U$$218/X sky130_fd_sc_hd__xor2_1
XFILLER_44_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater583 U$$1922/X VGND VGND VPWR VPWR U$$2046/A2 sky130_fd_sc_hd__buf_6
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$229 U$$92/A1 U$$263/A2 U$$94/A1 U$$231/B2 VGND VGND VPWR VPWR U$$230/A sky130_fd_sc_hd__a22o_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater594 U$$1746/A2 VGND VGND VPWR VPWR U$$1696/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_66_990 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_448 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1004 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_1192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1023 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1097 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_829 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_581 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_111_0 U$$3287/Y U$$3421/X U$$3554/X VGND VGND VPWR VPWR dadda_fa_4_112_1/A
+ dadda_fa_4_111_2/A sky130_fd_sc_hd__fa_1
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater1107 U$$3606/B1 VGND VGND VPWR VPWR U$$731/A1 sky130_fd_sc_hd__buf_8
Xrepeater1118 U$$44/A1 VGND VGND VPWR VPWR U$$866/A1 sky130_fd_sc_hd__buf_4
Xrepeater1129 input73/X VGND VGND VPWR VPWR U$$4289/A1 sky130_fd_sc_hd__buf_6
XFILLER_135_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_52_2 dadda_fa_3_52_2/A dadda_fa_3_52_2/B dadda_fa_3_52_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_1/A dadda_fa_4_52_2/B sky130_fd_sc_hd__fa_1
XFILLER_76_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_68_2 U$$1074/X U$$1207/X U$$1340/X VGND VGND VPWR VPWR dadda_fa_1_69_6/B
+ dadda_fa_1_68_8/A sky130_fd_sc_hd__fa_1
XTAP_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_45_1 dadda_fa_3_45_1/A dadda_fa_3_45_1/B dadda_fa_3_45_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_0/CIN dadda_fa_4_45_2/A sky130_fd_sc_hd__fa_1
XTAP_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_22_0 dadda_fa_6_22_0/A dadda_fa_6_22_0/B dadda_fa_6_22_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_23_0/B dadda_fa_7_22_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_60_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_38_0 dadda_fa_3_38_0/A dadda_fa_3_38_0/B dadda_fa_3_38_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_0/B dadda_fa_4_38_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$891 final_adder.U$$794/X final_adder.U$$503/X final_adder.U$$795/X
+ VGND VGND VPWR VPWR final_adder.U$$891/X sky130_fd_sc_hd__a21o_2
XU$$730 U$$730/A U$$750/B VGND VGND VPWR VPWR U$$730/X sky130_fd_sc_hd__xor2_1
XU$$741 U$$741/A1 U$$793/A2 U$$741/B1 U$$793/B2 VGND VGND VPWR VPWR U$$742/A sky130_fd_sc_hd__a22o_1
XFILLER_147_1210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$752 U$$752/A U$$796/B VGND VGND VPWR VPWR U$$752/X sky130_fd_sc_hd__xor2_1
XFILLER_17_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$763 U$$763/A1 U$$805/A2 U$$763/B1 U$$805/B2 VGND VGND VPWR VPWR U$$764/A sky130_fd_sc_hd__a22o_1
XFILLER_204_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$774 U$$774/A U$$794/B VGND VGND VPWR VPWR U$$774/X sky130_fd_sc_hd__xor2_1
XFILLER_32_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$785 U$$920/B1 U$$793/A2 U$$787/A1 U$$793/B2 VGND VGND VPWR VPWR U$$786/A sky130_fd_sc_hd__a22o_1
XU$$796 U$$796/A U$$796/B VGND VGND VPWR VPWR U$$796/X sky130_fd_sc_hd__xor2_1
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_176_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_2 _327_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdadda_fa_2_97_4 U$$3925/X U$$4058/X U$$4191/X VGND VGND VPWR VPWR dadda_fa_3_98_1/CIN
+ dadda_fa_3_97_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1630 U$$2206/B1 VGND VGND VPWR VPWR U$$975/A1 sky130_fd_sc_hd__buf_4
XFILLER_67_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1641 U$$2981/B1 VGND VGND VPWR VPWR U$$2159/B1 sky130_fd_sc_hd__buf_4
XFILLER_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1652 input107/X VGND VGND VPWR VPWR U$$4488/A1 sky130_fd_sc_hd__buf_4
Xrepeater1663 U$$4484/A1 VGND VGND VPWR VPWR U$$783/B1 sky130_fd_sc_hd__buf_4
XFILLER_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1674 U$$4480/B1 VGND VGND VPWR VPWR U$$3112/A1 sky130_fd_sc_hd__buf_6
XFILLER_153_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1685 U$$914/B1 VGND VGND VPWR VPWR U$$916/A1 sky130_fd_sc_hd__buf_6
XFILLER_28_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3979_1757 VGND VGND VPWR VPWR U$$3979_1757/HI U$$3979/A1 sky130_fd_sc_hd__conb_1
Xrepeater1696 U$$366/A1 VGND VGND VPWR VPWR U$$92/A1 sky130_fd_sc_hd__buf_4
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_40_0 U$$1550/X U$$1683/X U$$1816/X VGND VGND VPWR VPWR dadda_fa_3_41_0/B
+ dadda_fa_3_40_2/B sky130_fd_sc_hd__fa_1
XFILLER_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2170 U$$2170/A U$$2170/B VGND VGND VPWR VPWR U$$2170/X sky130_fd_sc_hd__xor2_1
XU$$2181 U$$4236/A1 U$$2183/A2 U$$4099/B1 U$$2183/B2 VGND VGND VPWR VPWR U$$2182/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2192 input25/X VGND VGND VPWR VPWR U$$2192/Y sky130_fd_sc_hd__inv_1
XFILLER_74_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1480 U$$930/B1 U$$1504/A2 U$$932/B1 U$$1504/B2 VGND VGND VPWR VPWR U$$1481/A sky130_fd_sc_hd__a22o_1
XU$$1491 U$$1491/A U$$1499/B VGND VGND VPWR VPWR U$$1491/X sky130_fd_sc_hd__xor2_1
XFILLER_210_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_2 U$$2305/X U$$2438/X U$$2571/X VGND VGND VPWR VPWR dadda_fa_2_86_3/A
+ dadda_fa_2_85_5/A sky130_fd_sc_hd__fa_1
XFILLER_104_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_62_1 dadda_fa_4_62_1/A dadda_fa_4_62_1/B dadda_fa_4_62_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/B dadda_fa_5_62_1/B sky130_fd_sc_hd__fa_1
Xdadda_fa_1_78_1 U$$1626/X U$$1759/X U$$1892/X VGND VGND VPWR VPWR dadda_fa_2_79_0/CIN
+ dadda_fa_2_78_3/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_4_55_0 dadda_fa_4_55_0/A dadda_fa_4_55_0/B dadda_fa_4_55_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/A dadda_fa_5_55_1/A sky130_fd_sc_hd__fa_1
XTAP_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$110 _406_/Q _278_/Q VGND VGND VPWR VPWR final_adder.U$$915/B1 final_adder.U$$144/A
+ sky130_fd_sc_hd__ha_1
XTAP_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$121 _417_/Q _289_/Q VGND VGND VPWR VPWR final_adder.U$$135/B1 final_adder.U$$134/B
+ sky130_fd_sc_hd__ha_2
XFILLER_100_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$132 final_adder.U$$132/A final_adder.U$$132/B VGND VGND VPWR VPWR
+ final_adder.U$$260/B sky130_fd_sc_hd__and2_1
XTAP_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$143 final_adder.U$$142/B final_adder.U$$913/B1 final_adder.U$$143/B1
+ VGND VGND VPWR VPWR final_adder.U$$143/X sky130_fd_sc_hd__a21o_1
XTAP_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$154 final_adder.U$$154/A final_adder.U$$154/B VGND VGND VPWR VPWR
+ final_adder.U$$282/B sky130_fd_sc_hd__and2_1
XTAP_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$165 final_adder.U$$164/B final_adder.U$$935/B1 final_adder.U$$165/B1
+ VGND VGND VPWR VPWR final_adder.U$$165/X sky130_fd_sc_hd__a21o_1
XTAP_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$176 final_adder.U$$176/A final_adder.U$$176/B VGND VGND VPWR VPWR
+ final_adder.U$$304/B sky130_fd_sc_hd__and2_1
XTAP_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$187 final_adder.U$$186/B final_adder.U$$957/B1 final_adder.U$$187/B1
+ VGND VGND VPWR VPWR final_adder.U$$187/X sky130_fd_sc_hd__a21o_1
XTAP_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1099 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater391 U$$1093/A2 VGND VGND VPWR VPWR U$$1083/A2 sky130_fd_sc_hd__buf_4
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$198 final_adder.U$$198/A final_adder.U$$198/B VGND VGND VPWR VPWR
+ final_adder.U$$326/B sky130_fd_sc_hd__and2_1
XTAP_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_382_ _382_/CLK _382_/D VGND VGND VPWR VPWR _382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_201_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_843 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _227_/CLK sky130_fd_sc_hd__clkbuf_8
Xdadda_ha_0_74_2 U$$1485/X U$$1618/X VGND VGND VPWR VPWR dadda_fa_1_75_8/B dadda_fa_2_74_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_108_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_73_0 U$$684/Y U$$818/X U$$951/X VGND VGND VPWR VPWR dadda_fa_1_74_7/B
+ dadda_fa_1_73_8/B sky130_fd_sc_hd__fa_1
XFILLER_0_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput150 c[119] VGND VGND VPWR VPWR input150/X sky130_fd_sc_hd__clkbuf_4
Xinput161 c[13] VGND VGND VPWR VPWR input161/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput172 c[23] VGND VGND VPWR VPWR input172/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput183 c[33] VGND VGND VPWR VPWR input183/X sky130_fd_sc_hd__clkbuf_4
XFILLER_209_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput194 c[43] VGND VGND VPWR VPWR input194/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1090 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$560 U$$969/B1 U$$578/A2 U$$836/A1 U$$578/B2 VGND VGND VPWR VPWR U$$561/A sky130_fd_sc_hd__a22o_1
XTAP_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$571 U$$571/A U$$607/B VGND VGND VPWR VPWR U$$571/X sky130_fd_sc_hd__xor2_1
XFILLER_17_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$582 U$$34/A1 U$$606/A2 U$$36/A1 U$$606/B2 VGND VGND VPWR VPWR U$$583/A sky130_fd_sc_hd__a22o_1
XU$$593 U$$593/A U$$625/B VGND VGND VPWR VPWR U$$593/X sky130_fd_sc_hd__xor2_1
XFILLER_204_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_665 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_692 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_95_1 U$$2990/X U$$3123/X U$$3256/X VGND VGND VPWR VPWR dadda_fa_3_96_0/CIN
+ dadda_fa_3_95_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_105_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_72_0 dadda_fa_5_72_0/A dadda_fa_5_72_0/B dadda_fa_5_72_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_73_0/A dadda_fa_6_72_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_2_88_0 U$$3508/X U$$3641/X U$$3774/X VGND VGND VPWR VPWR dadda_fa_3_89_0/B
+ dadda_fa_3_88_2/B sky130_fd_sc_hd__fa_1
XFILLER_67_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1460 U$$3451/A1 VGND VGND VPWR VPWR U$$2901/B1 sky130_fd_sc_hd__buf_4
XFILLER_132_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1471 U$$4408/A1 VGND VGND VPWR VPWR U$$4269/B1 sky130_fd_sc_hd__buf_6
XFILLER_160_559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1482 U$$4404/A1 VGND VGND VPWR VPWR U$$979/A1 sky130_fd_sc_hd__buf_4
Xrepeater1493 U$$3557/B1 VGND VGND VPWR VPWR U$$3283/B1 sky130_fd_sc_hd__buf_2
XFILLER_28_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_71_8 dadda_fa_1_71_8/A dadda_fa_1_71_8/B dadda_fa_1_71_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_72_3/A dadda_fa_3_71_0/A sky130_fd_sc_hd__fa_2
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_1028 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_7 dadda_fa_1_64_7/A dadda_fa_1_64_7/B dadda_fa_1_64_7/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_2/CIN dadda_fa_2_64_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_100_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_57_6 U$$3579/X U$$3712/X U$$3845/X VGND VGND VPWR VPWR dadda_fa_2_58_2/B
+ dadda_fa_2_57_5/B sky130_fd_sc_hd__fa_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_392 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_9_0 dadda_fa_7_9_0/A dadda_fa_7_9_0/B dadda_fa_7_9_0/CIN VGND VGND VPWR
+ VPWR _306_/D _177_/D sky130_fd_sc_hd__fa_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4244_1763 VGND VGND VPWR VPWR U$$4244_1763/HI U$$4244/B1 sky130_fd_sc_hd__conb_1
XFILLER_161_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_7_87_0 dadda_fa_7_87_0/A dadda_fa_7_87_0/B dadda_fa_7_87_0/CIN VGND VGND
+ VPWR VPWR _384_/D _255_/D sky130_fd_sc_hd__fa_2
XFILLER_136_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_90_0 dadda_fa_1_90_0/A U$$1916/X U$$2049/X VGND VGND VPWR VPWR dadda_fa_2_91_4/A
+ dadda_fa_2_90_5/A sky130_fd_sc_hd__fa_1
XFILLER_102_1190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_932 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4308 U$$4308/A U$$4382/B VGND VGND VPWR VPWR U$$4308/X sky130_fd_sc_hd__xor2_1
XU$$4319 U$$4456/A1 U$$4327/A2 U$$4458/A1 U$$4327/B2 VGND VGND VPWR VPWR U$$4320/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3607 U$$3607/A U$$3613/B VGND VGND VPWR VPWR U$$3607/X sky130_fd_sc_hd__xor2_1
XFILLER_46_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3618 input81/X U$$3660/A2 U$$3618/B1 U$$3660/B2 VGND VGND VPWR VPWR U$$3619/A
+ sky130_fd_sc_hd__a22o_1
XU$$3629 U$$3629/A input49/X VGND VGND VPWR VPWR U$$3629/X sky130_fd_sc_hd__xor2_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_6_102_0 dadda_fa_6_102_0/A dadda_fa_6_102_0/B dadda_fa_6_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_7_103_0/B dadda_fa_7_102_0/CIN sky130_fd_sc_hd__fa_1
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2906 U$$2906/A U$$2920/B VGND VGND VPWR VPWR U$$2906/X sky130_fd_sc_hd__xor2_1
XFILLER_46_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 _199_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2917 U$$4011/B1 U$$2919/A2 U$$4289/A1 U$$2919/B2 VGND VGND VPWR VPWR U$$2918/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2928 U$$2928/A U$$2950/B VGND VGND VPWR VPWR U$$2928/X sky130_fd_sc_hd__xor2_1
XANTENNA_211 _200_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2939 U$$3211/B1 U$$2967/A2 U$$3352/A1 U$$2967/B2 VGND VGND VPWR VPWR U$$2940/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_22_3 U$$1514/X U$$1574/B input171/X VGND VGND VPWR VPWR dadda_fa_4_23_1/B
+ dadda_fa_4_22_2/CIN sky130_fd_sc_hd__fa_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_244 _291_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 U$$4289/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_266 U$$3753/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_365_ _367_/CLK _365_/D VGND VGND VPWR VPWR _365_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_296_ _323_/CLK _296_/D VGND VGND VPWR VPWR _296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_67_5 dadda_fa_2_67_5/A dadda_fa_2_67_5/B dadda_fa_2_67_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_68_2/A dadda_fa_4_67_0/A sky130_fd_sc_hd__fa_2
XFILLER_84_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$390 U$$527/A1 U$$394/A2 U$$392/A1 U$$394/B2 VGND VGND VPWR VPWR U$$391/A sky130_fd_sc_hd__a22o_1
XFILLER_33_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1021 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1290 U$$3697/B VGND VGND VPWR VPWR U$$3623/B sky130_fd_sc_hd__buf_6
XFILLER_120_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_62_4 U$$3988/X U$$4121/X U$$4254/X VGND VGND VPWR VPWR dadda_fa_2_63_1/CIN
+ dadda_fa_2_62_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_55_3 U$$1979/X U$$2112/X U$$2245/X VGND VGND VPWR VPWR dadda_fa_2_56_1/B
+ dadda_fa_2_55_4/B sky130_fd_sc_hd__fa_1
XFILLER_132_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_690 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_32_2 dadda_fa_4_32_2/A dadda_fa_4_32_2/B dadda_fa_4_32_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_33_0/CIN dadda_fa_5_32_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_1_48_2 U$$901/X U$$1034/X U$$1167/X VGND VGND VPWR VPWR dadda_fa_2_49_1/CIN
+ dadda_fa_2_48_4/B sky130_fd_sc_hd__fa_1
XFILLER_82_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_25_1 dadda_fa_4_25_1/A dadda_fa_4_25_1/B dadda_fa_4_25_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/B dadda_fa_5_25_1/B sky130_fd_sc_hd__fa_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_18_0 U$$1107/X U$$1240/X U$$1272/B VGND VGND VPWR VPWR dadda_fa_5_19_0/A
+ dadda_fa_5_18_1/A sky130_fd_sc_hd__fa_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4105 U$$4379/A1 U$$4107/A2 U$$4242/B1 U$$4107/B2 VGND VGND VPWR VPWR U$$4106/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4116 U$$4116/A1 U$$4144/A2 U$$4392/A1 U$$4144/B2 VGND VGND VPWR VPWR U$$4117/A
+ sky130_fd_sc_hd__a22o_1
XU$$4127 U$$4127/A U$$4145/B VGND VGND VPWR VPWR U$$4127/X sky130_fd_sc_hd__xor2_1
XFILLER_24_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4138 U$$4275/A1 U$$4144/A2 U$$4275/B1 U$$4144/B2 VGND VGND VPWR VPWR U$$4139/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_150_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3404 input114/X U$$3422/A2 U$$3817/A1 U$$3422/B2 VGND VGND VPWR VPWR U$$3405/A
+ sky130_fd_sc_hd__a22o_1
XU$$4149 U$$4149/A U$$4189/B VGND VGND VPWR VPWR U$$4149/X sky130_fd_sc_hd__xor2_1
XU$$3415 U$$3415/A U$$3417/B VGND VGND VPWR VPWR U$$3415/X sky130_fd_sc_hd__xor2_1
XFILLER_58_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_392 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3426 input46/X VGND VGND VPWR VPWR U$$3428/B sky130_fd_sc_hd__inv_1
XFILLER_207_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3437 U$$3846/B1 U$$3527/A2 U$$3713/A1 U$$3527/B2 VGND VGND VPWR VPWR U$$3438/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2703 U$$2975/B1 U$$2607/X U$$2842/A1 U$$2608/X VGND VGND VPWR VPWR U$$2704/A sky130_fd_sc_hd__a22o_1
XFILLER_37_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3448 U$$3448/A U$$3454/B VGND VGND VPWR VPWR U$$3448/X sky130_fd_sc_hd__xor2_1
XU$$2714 U$$2714/A U$$2716/B VGND VGND VPWR VPWR U$$2714/X sky130_fd_sc_hd__xor2_1
XFILLER_37_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3459 U$$4005/B1 U$$3479/A2 U$$4009/A1 U$$3479/B2 VGND VGND VPWR VPWR U$$3460/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2725 U$$122/A1 U$$2735/A2 U$$3547/B1 U$$2735/B2 VGND VGND VPWR VPWR U$$2726/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2736 U$$2736/A U$$2736/B VGND VGND VPWR VPWR U$$2736/X sky130_fd_sc_hd__xor2_1
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2747 U$$2747/A U$$2755/B VGND VGND VPWR VPWR U$$2747/X sky130_fd_sc_hd__xor2_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2758 U$$3852/B1 U$$2790/A2 U$$3719/A1 U$$2790/B2 VGND VGND VPWR VPWR U$$2759/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_0 U$$47/X U$$180/X U$$313/X VGND VGND VPWR VPWR dadda_fa_4_21_0/B dadda_fa_4_20_1/CIN
+ sky130_fd_sc_hd__fa_1
XU$$2769 U$$2769/A U$$2783/B VGND VGND VPWR VPWR U$$2769/X sky130_fd_sc_hd__xor2_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1013 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_417_ _417_/CLK _417_/D VGND VGND VPWR VPWR _417_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_1185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_186_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_348_ _351_/CLK _348_/D VGND VGND VPWR VPWR _348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_1106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_279_ _408_/CLK _279_/D VGND VGND VPWR VPWR _279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_993 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_72_3 dadda_fa_2_72_3/A dadda_fa_2_72_3/B dadda_fa_2_72_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/B dadda_fa_3_72_3/B sky130_fd_sc_hd__fa_1
XFILLER_155_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_65_2 dadda_fa_2_65_2/A dadda_fa_2_65_2/B dadda_fa_2_65_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/A dadda_fa_3_65_3/A sky130_fd_sc_hd__fa_1
Xrepeater902 U$$4389/X VGND VGND VPWR VPWR U$$4512/B2 sky130_fd_sc_hd__buf_4
XFILLER_69_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$709 final_adder.U$$708/B final_adder.U$$605/X final_adder.U$$589/X
+ VGND VGND VPWR VPWR final_adder.U$$709/X sky130_fd_sc_hd__a21o_1
Xrepeater913 U$$3300/B1 VGND VGND VPWR VPWR U$$2069/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_42_1 dadda_fa_5_42_1/A dadda_fa_5_42_1/B dadda_fa_5_42_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_43_0/B dadda_fa_7_42_0/A sky130_fd_sc_hd__fa_2
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater924 U$$4468/B1 VGND VGND VPWR VPWR U$$3235/B1 sky130_fd_sc_hd__buf_6
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_2_58_1 dadda_fa_2_58_1/A dadda_fa_2_58_1/B dadda_fa_2_58_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_0/CIN dadda_fa_3_58_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater935 U$$4055/A1 VGND VGND VPWR VPWR U$$82/A1 sky130_fd_sc_hd__buf_6
Xrepeater946 U$$2957/A1 VGND VGND VPWR VPWR U$$3366/B1 sky130_fd_sc_hd__buf_8
XFILLER_110_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater957 U$$4049/B1 VGND VGND VPWR VPWR U$$3775/B1 sky130_fd_sc_hd__buf_4
Xrepeater968 U$$2951/A1 VGND VGND VPWR VPWR U$$483/B1 sky130_fd_sc_hd__buf_6
Xdadda_fa_5_35_0 dadda_fa_5_35_0/A dadda_fa_5_35_0/B dadda_fa_5_35_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_36_0/A dadda_fa_6_35_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_204_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater979 U$$4045/A1 VGND VGND VPWR VPWR U$$2810/B1 sky130_fd_sc_hd__buf_6
XFILLER_25_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3960 U$$3960/A1 U$$3966/A2 U$$3960/B1 U$$3966/B2 VGND VGND VPWR VPWR U$$3961/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3971 U$$3971/A U$$3971/B VGND VGND VPWR VPWR U$$3971/X sky130_fd_sc_hd__xor2_1
XFILLER_25_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2746_1738 VGND VGND VPWR VPWR U$$2746_1738/HI U$$2746/A1 sky130_fd_sc_hd__conb_1
XU$$3982 U$$3982/A U$$4012/B VGND VGND VPWR VPWR U$$3982/X sky130_fd_sc_hd__xor2_1
XU$$3993 U$$4402/B1 U$$4011/A2 U$$4269/A1 U$$4011/B2 VGND VGND VPWR VPWR U$$3994/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_180_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput262 output262/A VGND VGND VPWR VPWR o[104] sky130_fd_sc_hd__buf_2
Xdadda_fa_0_72_0_1849 VGND VGND VPWR VPWR dadda_fa_0_72_0/A dadda_fa_0_72_0_1849/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_88_911 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput273 output273/A VGND VGND VPWR VPWR o[114] sky130_fd_sc_hd__buf_2
XU$$3705_1753 VGND VGND VPWR VPWR U$$3705_1753/HI U$$3705/A1 sky130_fd_sc_hd__conb_1
Xoutput284 output284/A VGND VGND VPWR VPWR o[124] sky130_fd_sc_hd__buf_2
Xoutput295 output295/A VGND VGND VPWR VPWR o[19] sky130_fd_sc_hd__buf_2
XFILLER_82_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_60_1 U$$2388/X U$$2521/X U$$2654/X VGND VGND VPWR VPWR dadda_fa_2_61_0/CIN
+ dadda_fa_2_60_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_53_0 U$$379/X U$$512/X U$$645/X VGND VGND VPWR VPWR dadda_fa_2_54_0/B
+ dadda_fa_2_53_3/B sky130_fd_sc_hd__fa_1
XFILLER_56_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1309 U$$1446/A1 U$$1311/A2 U$$1448/A1 U$$1355/B2 VGND VGND VPWR VPWR U$$1310/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1024_1846 VGND VGND VPWR VPWR final_adder.U$$1024_1846/HI final_adder.U$$1024/B
+ sky130_fd_sc_hd__conb_1
XFILLER_128_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_202_ _337_/CLK _202_/D VGND VGND VPWR VPWR _202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1103 final_adder.U$$176/B final_adder.U$$947/X VGND VGND VPWR VPWR
+ output361/A sky130_fd_sc_hd__xor2_1
XFILLER_183_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$1114 final_adder.U$$164/A ANTENNA_250/DIODE VGND VGND VPWR VPWR output374/A
+ sky130_fd_sc_hd__xor2_1
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1125 final_adder.U$$154/B final_adder.U$$925/X VGND VGND VPWR VPWR
+ output259/A sky130_fd_sc_hd__xor2_2
Xfinal_adder.U$$1136 final_adder.U$$142/A final_adder.U$$851/X VGND VGND VPWR VPWR
+ output271/A sky130_fd_sc_hd__xor2_1
XFILLER_184_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1147 final_adder.U$$132/B final_adder.U$$903/X VGND VGND VPWR VPWR
+ output283/A sky130_fd_sc_hd__xor2_1
XFILLER_165_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_695 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_82_2 dadda_fa_3_82_2/A dadda_fa_3_82_2/B dadda_fa_3_82_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_1/A dadda_fa_4_82_2/B sky130_fd_sc_hd__fa_1
XFILLER_48_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_75_1 dadda_fa_3_75_1/A dadda_fa_3_75_1/B dadda_fa_3_75_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_0/CIN dadda_fa_4_75_2/A sky130_fd_sc_hd__fa_1
XFILLER_174_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_52_0 dadda_fa_6_52_0/A dadda_fa_6_52_0/B dadda_fa_6_52_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_53_0/B dadda_fa_7_52_0/CIN sky130_fd_sc_hd__fa_2
Xdadda_fa_3_68_0 dadda_fa_3_68_0/A dadda_fa_3_68_0/B dadda_fa_3_68_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_0/B dadda_fa_4_68_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_61_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3201 U$$4434/A1 U$$3207/A2 U$$4297/B1 U$$3207/B2 VGND VGND VPWR VPWR U$$3202/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$3212 U$$3212/A U$$3228/B VGND VGND VPWR VPWR U$$3212/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_4_111_2 dadda_fa_4_111_2/A dadda_fa_4_111_2/B dadda_fa_4_111_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_112_0/CIN dadda_fa_5_111_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_150_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3223 U$$4045/A1 U$$3155/X input91/X U$$3156/X VGND VGND VPWR VPWR U$$3224/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$16 _312_/Q _184_/Q VGND VGND VPWR VPWR final_adder.U$$239/A2 final_adder.U$$238/A
+ sky130_fd_sc_hd__ha_1
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3234 U$$3234/A U$$3242/B VGND VGND VPWR VPWR U$$3234/X sky130_fd_sc_hd__xor2_1
XFILLER_206_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2500 U$$3183/B1 U$$2596/A2 U$$719/B1 U$$2596/B2 VGND VGND VPWR VPWR U$$2501/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3245 U$$3245/A1 U$$3155/X U$$3245/B1 U$$3156/X VGND VGND VPWR VPWR U$$3246/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$27 _323_/Q _195_/Q VGND VGND VPWR VPWR final_adder.U$$229/B1 final_adder.U$$228/B
+ sky130_fd_sc_hd__ha_1
XU$$3256 U$$3256/A U$$3256/B VGND VGND VPWR VPWR U$$3256/X sky130_fd_sc_hd__xor2_1
XU$$2511 U$$2511/A U$$2597/B VGND VGND VPWR VPWR U$$2511/X sky130_fd_sc_hd__xor2_1
XFILLER_98_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_104_1 dadda_fa_4_104_1/A dadda_fa_4_104_1/B dadda_fa_4_104_1/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/B dadda_fa_5_104_1/B sky130_fd_sc_hd__fa_1
XU$$3267 U$$116/A1 U$$3285/A2 U$$3680/A1 U$$3285/B2 VGND VGND VPWR VPWR U$$3268/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$38 _334_/Q _206_/Q VGND VGND VPWR VPWR final_adder.U$$987/B1 final_adder.U$$216/A
+ sky130_fd_sc_hd__ha_1
XU$$2522 U$$330/A1 U$$2542/A2 U$$3207/B1 U$$2542/B2 VGND VGND VPWR VPWR U$$2523/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$49 _345_/Q _217_/Q VGND VGND VPWR VPWR final_adder.U$$207/B1 final_adder.U$$206/B
+ sky130_fd_sc_hd__ha_1
XU$$2533 U$$2533/A U$$2577/B VGND VGND VPWR VPWR U$$2533/X sky130_fd_sc_hd__xor2_1
XFILLER_46_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3278 U$$3278/A U$$3287/A VGND VGND VPWR VPWR U$$3278/X sky130_fd_sc_hd__xor2_1
XFILLER_206_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2544 U$$2955/A1 U$$2558/A2 U$$2957/A1 U$$2558/B2 VGND VGND VPWR VPWR U$$2545/A
+ sky130_fd_sc_hd__a22o_1
XU$$3289 input43/X VGND VGND VPWR VPWR U$$3291/B sky130_fd_sc_hd__inv_1
XFILLER_94_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2555 U$$2555/A U$$2601/B VGND VGND VPWR VPWR U$$2555/X sky130_fd_sc_hd__xor2_1
XU$$1810 U$$1810/A U$$1832/B VGND VGND VPWR VPWR U$$1810/X sky130_fd_sc_hd__xor2_1
XU$$1821 U$$860/B1 U$$1869/A2 U$$727/A1 U$$1869/B2 VGND VGND VPWR VPWR U$$1822/A sky130_fd_sc_hd__a22o_1
XU$$2566 U$$3114/A1 U$$2470/X U$$3116/A1 U$$2471/X VGND VGND VPWR VPWR U$$2567/A sky130_fd_sc_hd__a22o_1
XU$$2577 U$$2577/A U$$2577/B VGND VGND VPWR VPWR U$$2577/X sky130_fd_sc_hd__xor2_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1832 U$$1832/A U$$1832/B VGND VGND VPWR VPWR U$$1832/X sky130_fd_sc_hd__xor2_1
XU$$2588 U$$4095/A1 U$$2588/A2 U$$3960/A1 U$$2588/B2 VGND VGND VPWR VPWR U$$2589/A
+ sky130_fd_sc_hd__a22o_1
XU$$1843 U$$3348/B1 U$$1879/A2 U$$3215/A1 U$$1879/B2 VGND VGND VPWR VPWR U$$1844/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1854 U$$1854/A U$$1880/B VGND VGND VPWR VPWR U$$1854/X sky130_fd_sc_hd__xor2_1
XFILLER_210_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2599 U$$2599/A U$$2601/B VGND VGND VPWR VPWR U$$2599/X sky130_fd_sc_hd__xor2_1
XFILLER_15_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$1865 U$$3235/A1 U$$1785/X U$$3235/B1 U$$1786/X VGND VGND VPWR VPWR U$$1866/A sky130_fd_sc_hd__a22o_1
XU$$1876 U$$1876/A U$$1878/B VGND VGND VPWR VPWR U$$1876/X sky130_fd_sc_hd__xor2_1
XU$$1887 U$$517/A1 U$$1915/A2 U$$517/B1 U$$1915/B2 VGND VGND VPWR VPWR U$$1888/A sky130_fd_sc_hd__a22o_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1898 U$$1898/A U$$1917/A VGND VGND VPWR VPWR U$$1898/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_7_125_0 dadda_fa_7_125_0/A dadda_fa_7_125_0/B dadda_fa_7_125_0/CIN VGND
+ VGND VPWR VPWR _422_/D _293_/D sky130_fd_sc_hd__fa_1
XFILLER_203_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_70_0 dadda_fa_2_70_0/A dadda_fa_2_70_0/B dadda_fa_2_70_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_0/B dadda_fa_3_70_2/B sky130_fd_sc_hd__fa_1
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater710 U$$3753/B2 VGND VGND VPWR VPWR U$$3793/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$517 final_adder.U$$516/B final_adder.U$$401/X final_adder.U$$393/X
+ VGND VGND VPWR VPWR final_adder.U$$517/X sky130_fd_sc_hd__a21o_1
Xrepeater721 U$$3686/B2 VGND VGND VPWR VPWR U$$3680/B2 sky130_fd_sc_hd__buf_4
XFILLER_69_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$528 final_adder.U$$536/B final_adder.U$$528/B VGND VGND VPWR VPWR
+ final_adder.U$$648/B sky130_fd_sc_hd__and2_1
Xrepeater732 U$$3517/B2 VGND VGND VPWR VPWR U$$3489/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$539 final_adder.U$$538/B final_adder.U$$423/X final_adder.U$$415/X
+ VGND VGND VPWR VPWR final_adder.U$$539/X sky130_fd_sc_hd__a21o_1
Xrepeater743 U$$3241/B2 VGND VGND VPWR VPWR U$$3207/B2 sky130_fd_sc_hd__buf_12
Xrepeater754 U$$3132/B2 VGND VGND VPWR VPWR U$$3148/B2 sky130_fd_sc_hd__buf_6
Xrepeater765 U$$2882/X VGND VGND VPWR VPWR U$$2985/B2 sky130_fd_sc_hd__buf_6
Xrepeater776 U$$2844/B2 VGND VGND VPWR VPWR U$$2810/B2 sky130_fd_sc_hd__buf_6
XFILLER_84_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater787 U$$2735/B2 VGND VGND VPWR VPWR U$$2727/B2 sky130_fd_sc_hd__buf_6
XFILLER_72_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$4480 input103/X U$$4388/X U$$4480/B1 U$$4486/B2 VGND VGND VPWR VPWR U$$4481/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater798 U$$2471/X VGND VGND VPWR VPWR U$$2576/B2 sky130_fd_sc_hd__buf_6
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4491 U$$4491/A U$$4491/B VGND VGND VPWR VPWR U$$4491/X sky130_fd_sc_hd__xor2_1
XFILLER_71_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3790 U$$3790/A U$$3794/B VGND VGND VPWR VPWR U$$3790/X sky130_fd_sc_hd__xor2_1
XFILLER_53_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_674 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_359 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_166_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1025 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_92_1 dadda_fa_4_92_1/A dadda_fa_4_92_1/B dadda_fa_4_92_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/B dadda_fa_5_92_1/B sky130_fd_sc_hd__fa_1
XFILLER_10_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_610 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_85_0 dadda_fa_4_85_0/A dadda_fa_4_85_0/B dadda_fa_4_85_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/A dadda_fa_5_85_1/A sky130_fd_sc_hd__fa_1
XFILLER_109_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_106_3 dadda_fa_3_106_3/A dadda_fa_3_106_3/B dadda_fa_3_106_3/CIN VGND
+ VGND VPWR VPWR dadda_fa_4_107_1/B dadda_fa_4_106_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_107_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_161_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$901 U$$901/A U$$951/B VGND VGND VPWR VPWR U$$901/X sky130_fd_sc_hd__xor2_1
XU$$912 U$$912/A1 U$$918/A2 U$$914/A1 U$$918/B2 VGND VGND VPWR VPWR U$$913/A sky130_fd_sc_hd__a22o_1
XU$$923 U$$923/A U$$951/B VGND VGND VPWR VPWR U$$923/X sky130_fd_sc_hd__xor2_1
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$934 U$$934/A1 U$$826/X U$$936/A1 U$$827/X VGND VGND VPWR VPWR U$$935/A sky130_fd_sc_hd__a22o_1
XU$$945 U$$945/A U$$945/B VGND VGND VPWR VPWR U$$945/X sky130_fd_sc_hd__xor2_1
XFILLER_43_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$956 U$$956/A1 U$$826/X U$$956/B1 U$$827/X VGND VGND VPWR VPWR U$$957/A sky130_fd_sc_hd__a22o_1
XFILLER_204_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$967 U$$967/A1 U$$979/A2 U$$969/A1 U$$979/B2 VGND VGND VPWR VPWR U$$968/A sky130_fd_sc_hd__a22o_1
XU$$1106 U$$8/B1 U$$1138/A2 U$$12/A1 U$$1138/B2 VGND VGND VPWR VPWR U$$1107/A sky130_fd_sc_hd__a22o_1
XFILLER_189_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1117 U$$1117/A U$$1137/B VGND VGND VPWR VPWR U$$1117/X sky130_fd_sc_hd__xor2_1
XU$$978 U$$978/A U$$980/B VGND VGND VPWR VPWR U$$978/X sky130_fd_sc_hd__xor2_1
XFILLER_203_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1128 U$$991/A1 U$$1136/A2 U$$2363/A1 U$$1136/B2 VGND VGND VPWR VPWR U$$1129/A
+ sky130_fd_sc_hd__a22o_1
XU$$989 U$$989/A1 U$$993/A2 U$$991/A1 U$$993/B2 VGND VGND VPWR VPWR U$$990/A sky130_fd_sc_hd__a22o_1
XFILLER_189_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1139 U$$1139/A U$$1139/B VGND VGND VPWR VPWR U$$1139/X sky130_fd_sc_hd__xor2_1
XFILLER_43_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_188_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1081 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_882 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_169_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_996 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_860 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_42_4 dadda_fa_2_42_4/A dadda_fa_2_42_4/B dadda_fa_2_42_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_43_1/CIN dadda_fa_3_42_3/CIN sky130_fd_sc_hd__fa_1
XU$$3020 U$$3020/A1 U$$3060/A2 U$$3159/A1 U$$3060/B2 VGND VGND VPWR VPWR U$$3021/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$3031 U$$3031/A U$$3083/B VGND VGND VPWR VPWR U$$3031/X sky130_fd_sc_hd__xor2_1
XFILLER_207_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3042 input66/X U$$3124/A2 U$$30/A1 U$$3124/B2 VGND VGND VPWR VPWR U$$3043/A sky130_fd_sc_hd__a22o_1
XFILLER_53_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3053 U$$3053/A U$$3083/B VGND VGND VPWR VPWR U$$3053/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_35_3 U$$1540/X U$$1673/X U$$1806/X VGND VGND VPWR VPWR dadda_fa_3_36_1/B
+ dadda_fa_3_35_3/B sky130_fd_sc_hd__fa_1
XU$$3064 U$$4434/A1 U$$3108/A2 U$$4436/A1 U$$3108/B2 VGND VGND VPWR VPWR U$$3065/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$2330 input28/X VGND VGND VPWR VPWR U$$2332/B sky130_fd_sc_hd__inv_1
XU$$3075 U$$3075/A U$$3075/B VGND VGND VPWR VPWR U$$3075/X sky130_fd_sc_hd__xor2_1
XFILLER_207_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3086 U$$4456/A1 U$$3118/A2 U$$3088/A1 U$$3118/B2 VGND VGND VPWR VPWR U$$3087/A
+ sky130_fd_sc_hd__a22o_1
XU$$2341 U$$3300/A1 U$$2359/A2 U$$3300/B1 U$$2359/B2 VGND VGND VPWR VPWR U$$2342/A
+ sky130_fd_sc_hd__a22o_1
XU$$2352 U$$2352/A U$$2360/B VGND VGND VPWR VPWR U$$2352/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_28_2 U$$861/X U$$994/X U$$1127/X VGND VGND VPWR VPWR dadda_fa_3_29_2/B
+ dadda_fa_3_28_3/CIN sky130_fd_sc_hd__fa_1
XU$$3097 U$$3097/A U$$3151/A VGND VGND VPWR VPWR U$$3097/X sky130_fd_sc_hd__xor2_1
XU$$2363 U$$2363/A1 U$$2417/A2 U$$995/A1 U$$2417/B2 VGND VGND VPWR VPWR U$$2364/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2374 U$$2374/A U$$2380/B VGND VGND VPWR VPWR U$$2374/X sky130_fd_sc_hd__xor2_1
XFILLER_34_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1640 U$$1640/A U$$1644/A VGND VGND VPWR VPWR U$$1640/X sky130_fd_sc_hd__xor2_1
XFILLER_50_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2385 U$$741/A1 U$$2417/A2 U$$741/B1 U$$2417/B2 VGND VGND VPWR VPWR U$$2386/A sky130_fd_sc_hd__a22o_1
XU$$2396 U$$2396/A U$$2442/B VGND VGND VPWR VPWR U$$2396/X sky130_fd_sc_hd__xor2_1
XU$$1651 U$$1651/A U$$1679/B VGND VGND VPWR VPWR U$$1651/X sky130_fd_sc_hd__xor2_1
XU$$4381_1765 VGND VGND VPWR VPWR U$$4381_1765/HI U$$4381/B1 sky130_fd_sc_hd__conb_1
XU$$1662 U$$1799/A1 U$$1696/A2 U$$1799/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1663/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1673 U$$1673/A U$$1707/B VGND VGND VPWR VPWR U$$1673/X sky130_fd_sc_hd__xor2_1
XFILLER_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1684 U$$860/B1 U$$1688/A2 U$$727/A1 U$$1688/B2 VGND VGND VPWR VPWR U$$1685/A sky130_fd_sc_hd__a22o_1
XFILLER_148_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1695 U$$1695/A U$$1751/B VGND VGND VPWR VPWR U$$1695/X sky130_fd_sc_hd__xor2_1
XFILLER_124_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_187_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$303 final_adder.U$$302/B final_adder.U$$177/X final_adder.U$$175/X
+ VGND VGND VPWR VPWR final_adder.U$$303/X sky130_fd_sc_hd__a21o_1
XTAP_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$314 final_adder.U$$316/B final_adder.U$$314/B VGND VGND VPWR VPWR
+ final_adder.U$$440/B sky130_fd_sc_hd__and2_1
XFILLER_131_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$325 final_adder.U$$324/B final_adder.U$$199/X final_adder.U$$197/X
+ VGND VGND VPWR VPWR final_adder.U$$325/X sky130_fd_sc_hd__a21o_1
XFILLER_58_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$336 final_adder.U$$338/B final_adder.U$$336/B VGND VGND VPWR VPWR
+ final_adder.U$$462/B sky130_fd_sc_hd__and2_1
Xrepeater540 U$$2735/A2 VGND VGND VPWR VPWR U$$2727/A2 sky130_fd_sc_hd__buf_6
XTAP_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$347 final_adder.U$$346/B final_adder.U$$221/X final_adder.U$$219/X
+ VGND VGND VPWR VPWR final_adder.U$$347/X sky130_fd_sc_hd__a21o_1
XTAP_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater551 U$$2470/X VGND VGND VPWR VPWR U$$2576/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$358 final_adder.U$$360/B final_adder.U$$358/B VGND VGND VPWR VPWR
+ final_adder.U$$484/B sky130_fd_sc_hd__and2_1
XTAP_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater562 U$$2302/A2 VGND VGND VPWR VPWR U$$2272/A2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$369 final_adder.U$$368/B final_adder.U$$243/X final_adder.U$$241/X
+ VGND VGND VPWR VPWR final_adder.U$$369/X sky130_fd_sc_hd__a21o_1
Xrepeater573 U$$2059/X VGND VGND VPWR VPWR U$$2183/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_84_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$208 U$$208/A U$$212/B VGND VGND VPWR VPWR U$$208/X sky130_fd_sc_hd__xor2_1
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater584 U$$1869/A2 VGND VGND VPWR VPWR U$$1819/A2 sky130_fd_sc_hd__buf_4
XU$$219 U$$630/A1 U$$263/A2 U$$630/B1 U$$231/B2 VGND VGND VPWR VPWR U$$220/A sky130_fd_sc_hd__a22o_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater595 U$$1750/A2 VGND VGND VPWR VPWR U$$1706/A2 sky130_fd_sc_hd__buf_6
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1016 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_164_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1108 input75/X VGND VGND VPWR VPWR U$$3606/B1 sky130_fd_sc_hd__clkbuf_8
Xdadda_fa_3_111_1 U$$3687/X U$$3820/X U$$3953/X VGND VGND VPWR VPWR dadda_fa_4_112_1/B
+ dadda_fa_4_111_2/B sky130_fd_sc_hd__fa_1
XFILLER_112_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1119 U$$4015/B1 VGND VGND VPWR VPWR U$$44/A1 sky130_fd_sc_hd__buf_6
XFILLER_14_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_104_0 U$$3806/X U$$3939/X U$$4072/X VGND VGND VPWR VPWR dadda_fa_4_105_0/B
+ dadda_fa_4_104_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_88_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1058 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_56 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_3_52_3 dadda_fa_3_52_3/A dadda_fa_3_52_3/B dadda_fa_3_52_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_53_1/B dadda_fa_4_52_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_0_68_3 U$$1473/X U$$1606/X U$$1739/X VGND VGND VPWR VPWR dadda_fa_1_69_6/CIN
+ dadda_fa_1_68_8/B sky130_fd_sc_hd__fa_1
XFILLER_76_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_45_2 dadda_fa_3_45_2/A dadda_fa_3_45_2/B dadda_fa_3_45_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_1/A dadda_fa_4_45_2/B sky130_fd_sc_hd__fa_1
XFILLER_75_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$881 final_adder.U$$784/X final_adder.U$$737/X final_adder.U$$785/X
+ VGND VGND VPWR VPWR final_adder.U$$881/X sky130_fd_sc_hd__a21o_2
Xdadda_fa_3_38_1 dadda_fa_3_38_1/A dadda_fa_3_38_1/B dadda_fa_3_38_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_0/CIN dadda_fa_4_38_2/A sky130_fd_sc_hd__fa_1
XU$$720 U$$720/A U$$740/B VGND VGND VPWR VPWR U$$720/X sky130_fd_sc_hd__xor2_1
XU$$731 U$$731/A1 U$$739/A2 U$$733/A1 U$$739/B2 VGND VGND VPWR VPWR U$$732/A sky130_fd_sc_hd__a22o_1
XFILLER_95_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$742 U$$742/A U$$770/B VGND VGND VPWR VPWR U$$742/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_6_15_0 dadda_fa_6_15_0/A dadda_fa_6_15_0/B dadda_fa_6_15_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_16_0/B dadda_fa_7_15_0/CIN sky130_fd_sc_hd__fa_1
Xclkbuf_leaf_55_clk clkbuf_3_1_0_clk/X VGND VGND VPWR VPWR _362_/CLK sky130_fd_sc_hd__clkbuf_16
XU$$753 U$$890/A1 U$$759/A2 U$$892/A1 U$$759/B2 VGND VGND VPWR VPWR U$$754/A sky130_fd_sc_hd__a22o_1
XFILLER_182_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$764 U$$764/A U$$796/B VGND VGND VPWR VPWR U$$764/X sky130_fd_sc_hd__xor2_1
XFILLER_72_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$775 U$$912/A1 U$$783/A2 U$$914/A1 U$$783/B2 VGND VGND VPWR VPWR U$$776/A sky130_fd_sc_hd__a22o_1
XFILLER_147_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$786 U$$786/A U$$794/B VGND VGND VPWR VPWR U$$786/X sky130_fd_sc_hd__xor2_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$797 U$$932/B1 U$$805/A2 U$$799/A1 U$$805/B2 VGND VGND VPWR VPWR U$$798/A sky130_fd_sc_hd__a22o_1
XFILLER_32_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_1029 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_ha_3_110_3 U$$4350/X U$$4483/X VGND VGND VPWR VPWR dadda_fa_4_111_1/CIN dadda_ha_3_110_3/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_32_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_499 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_177_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_3 _327_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_2_97_5 U$$4324/X U$$4457/X input253/X VGND VGND VPWR VPWR dadda_fa_3_98_2/A
+ dadda_fa_4_97_0/A sky130_fd_sc_hd__fa_2
Xrepeater1620 U$$1286/B VGND VGND VPWR VPWR U$$1270/B sky130_fd_sc_hd__buf_6
XFILLER_160_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1631 input109/X VGND VGND VPWR VPWR U$$2206/B1 sky130_fd_sc_hd__buf_4
XFILLER_193_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_160_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1642 U$$4490/A1 VGND VGND VPWR VPWR U$$2981/B1 sky130_fd_sc_hd__buf_4
Xrepeater1653 U$$4484/B1 VGND VGND VPWR VPWR U$$4210/B1 sky130_fd_sc_hd__buf_4
XFILLER_153_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1664 U$$2701/B1 VGND VGND VPWR VPWR U$$98/B1 sky130_fd_sc_hd__buf_6
Xrepeater1675 U$$4480/B1 VGND VGND VPWR VPWR U$$783/A1 sky130_fd_sc_hd__buf_8
XFILLER_113_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater1686 U$$4478/A1 VGND VGND VPWR VPWR U$$914/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1697 U$$366/A1 VGND VGND VPWR VPWR U$$2967/B1 sky130_fd_sc_hd__buf_8
XFILLER_154_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_40_1 U$$1949/X U$$2082/X U$$2215/X VGND VGND VPWR VPWR dadda_fa_3_41_0/CIN
+ dadda_fa_3_40_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_33_0 U$$73/X U$$206/X U$$339/X VGND VGND VPWR VPWR dadda_fa_3_34_0/B dadda_fa_3_33_2/B
+ sky130_fd_sc_hd__fa_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2160 U$$2160/A U$$2184/B VGND VGND VPWR VPWR U$$2160/X sky130_fd_sc_hd__xor2_1
XU$$2171 U$$936/B1 U$$2177/A2 U$$2445/B1 U$$2177/B2 VGND VGND VPWR VPWR U$$2172/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2182 U$$2182/A U$$2184/B VGND VGND VPWR VPWR U$$2182/X sky130_fd_sc_hd__xor2_1
XU$$2193 input26/X VGND VGND VPWR VPWR U$$2195/B sky130_fd_sc_hd__inv_1
XU$$1470 U$$2975/B1 U$$1470/A2 U$$2842/A1 U$$1470/B2 VGND VGND VPWR VPWR U$$1471/A
+ sky130_fd_sc_hd__a22o_1
XU$$1481 U$$1481/A U$$1501/B VGND VGND VPWR VPWR U$$1481/X sky130_fd_sc_hd__xor2_1
XFILLER_50_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1492 U$$1764/B1 U$$1502/A2 U$$946/A1 U$$1502/B2 VGND VGND VPWR VPWR U$$1493/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_ha_1_86_5 U$$3504/X U$$3637/X VGND VGND VPWR VPWR dadda_fa_2_87_4/B dadda_fa_3_86_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_176_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$1513_1719 VGND VGND VPWR VPWR U$$1513_1719/HI U$$1513/A1 sky130_fd_sc_hd__conb_1
XFILLER_191_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_933 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_171_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_3 U$$2704/X U$$2837/X U$$2970/X VGND VGND VPWR VPWR dadda_fa_2_86_3/B
+ dadda_fa_2_85_5/B sky130_fd_sc_hd__fa_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_62_2 dadda_fa_4_62_2/A dadda_fa_4_62_2/B dadda_fa_4_62_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_63_0/CIN dadda_fa_5_62_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_89_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_1_78_2 U$$2025/X U$$2158/X U$$2291/X VGND VGND VPWR VPWR dadda_fa_2_79_1/A
+ dadda_fa_2_78_4/A sky130_fd_sc_hd__fa_1
XFILLER_103_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_55_1 dadda_fa_4_55_1/A dadda_fa_4_55_1/B dadda_fa_4_55_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/B dadda_fa_5_55_1/B sky130_fd_sc_hd__fa_1
XTAP_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfinal_adder.U$$100 _396_/Q _268_/Q VGND VGND VPWR VPWR final_adder.U$$925/B1 final_adder.U$$154/A
+ sky130_fd_sc_hd__ha_1
XTAP_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$111 _407_/Q _279_/Q VGND VGND VPWR VPWR final_adder.U$$145/B1 final_adder.U$$144/B
+ sky130_fd_sc_hd__ha_1
XTAP_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_32_0 dadda_fa_7_32_0/A dadda_fa_7_32_0/B dadda_fa_7_32_0/CIN VGND VGND
+ VPWR VPWR _329_/D _200_/D sky130_fd_sc_hd__fa_2
XFILLER_170_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$122 _418_/Q _290_/Q VGND VGND VPWR VPWR final_adder.U$$903/B1 final_adder.U$$132/A
+ sky130_fd_sc_hd__ha_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_48_0 dadda_fa_4_48_0/A dadda_fa_4_48_0/B dadda_fa_4_48_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/A dadda_fa_5_48_1/A sky130_fd_sc_hd__fa_1
Xfinal_adder.U$$133 final_adder.U$$132/B final_adder.U$$903/B1 final_adder.U$$133/B1
+ VGND VGND VPWR VPWR final_adder.U$$133/X sky130_fd_sc_hd__a21o_1
XTAP_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$144 final_adder.U$$144/A final_adder.U$$144/B VGND VGND VPWR VPWR
+ final_adder.U$$272/B sky130_fd_sc_hd__and2_1
XTAP_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$155 final_adder.U$$154/B final_adder.U$$925/B1 final_adder.U$$155/B1
+ VGND VGND VPWR VPWR final_adder.U$$155/X sky130_fd_sc_hd__a21o_1
XTAP_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$166 final_adder.U$$166/A final_adder.U$$166/B VGND VGND VPWR VPWR
+ final_adder.U$$294/B sky130_fd_sc_hd__and2_1
XTAP_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$177 final_adder.U$$176/B final_adder.U$$947/B1 final_adder.U$$177/B1
+ VGND VGND VPWR VPWR final_adder.U$$177/X sky130_fd_sc_hd__a21o_1
XTAP_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$188 final_adder.U$$188/A final_adder.U$$188/B VGND VGND VPWR VPWR
+ final_adder.U$$316/B sky130_fd_sc_hd__and2_1
XTAP_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater392 U$$963/X VGND VGND VPWR VPWR U$$1093/A2 sky130_fd_sc_hd__buf_8
XFILLER_211_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$199 final_adder.U$$198/B final_adder.U$$969/B1 final_adder.U$$199/B1
+ VGND VGND VPWR VPWR final_adder.U$$199/X sky130_fd_sc_hd__a21o_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_37_clk _239_/CLK VGND VGND VPWR VPWR _377_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_381_ _381_/CLK _381_/D VGND VGND VPWR VPWR _381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_182_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_120_0_1869 VGND VGND VPWR VPWR dadda_fa_4_120_0/A dadda_fa_4_120_0_1869/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_141_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_0_73_1 U$$1084/X U$$1217/X U$$1350/X VGND VGND VPWR VPWR dadda_fa_1_74_7/CIN
+ dadda_fa_1_73_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_209_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput140 c[10] VGND VGND VPWR VPWR input140/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_3_50_0 dadda_fa_3_50_0/A dadda_fa_3_50_0/B dadda_fa_3_50_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_0/B dadda_fa_4_50_1/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_0_66_0 U$$136/A U$$272/X U$$405/X VGND VGND VPWR VPWR dadda_fa_1_67_5/B
+ dadda_fa_1_66_7/B sky130_fd_sc_hd__fa_1
XFILLER_23_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput151 c[11] VGND VGND VPWR VPWR input151/X sky130_fd_sc_hd__clkbuf_4
Xinput162 c[14] VGND VGND VPWR VPWR input162/X sky130_fd_sc_hd__clkbuf_4
Xinput173 c[24] VGND VGND VPWR VPWR input173/X sky130_fd_sc_hd__buf_2
XTAP_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput184 c[34] VGND VGND VPWR VPWR input184/X sky130_fd_sc_hd__buf_2
XTAP_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput195 c[44] VGND VGND VPWR VPWR input195/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_clk _255_/CLK VGND VGND VPWR VPWR _411_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$550 U$$685/A VGND VGND VPWR VPWR U$$550/Y sky130_fd_sc_hd__inv_1
XFILLER_45_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$561 U$$561/A U$$579/B VGND VGND VPWR VPWR U$$561/X sky130_fd_sc_hd__xor2_1
XTAP_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$572 U$$983/A1 U$$606/A2 U$$846/B1 U$$606/B2 VGND VGND VPWR VPWR U$$573/A sky130_fd_sc_hd__a22o_1
XFILLER_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$583 U$$583/A U$$607/B VGND VGND VPWR VPWR U$$583/X sky130_fd_sc_hd__xor2_1
XU$$594 U$$594/A1 U$$624/A2 U$$594/B1 U$$624/B2 VGND VGND VPWR VPWR U$$595/A sky130_fd_sc_hd__a22o_1
XFILLER_72_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_677 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_1214 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_95_2 U$$3389/X U$$3522/X U$$3655/X VGND VGND VPWR VPWR dadda_fa_3_96_1/A
+ dadda_fa_3_95_3/A sky130_fd_sc_hd__fa_1
XFILLER_145_579 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3842_1755 VGND VGND VPWR VPWR U$$3842_1755/HI U$$3842/A1 sky130_fd_sc_hd__conb_1
Xrepeater1450 U$$1507/A VGND VGND VPWR VPWR U$$1506/A sky130_fd_sc_hd__buf_8
Xdadda_fa_5_72_1 dadda_fa_5_72_1/A dadda_fa_5_72_1/B dadda_fa_5_72_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_73_0/B dadda_fa_7_72_0/A sky130_fd_sc_hd__fa_1
Xrepeater1461 U$$3451/A1 VGND VGND VPWR VPWR U$$26/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_88_1 U$$3907/X U$$4040/X U$$4173/X VGND VGND VPWR VPWR dadda_fa_3_89_0/CIN
+ dadda_fa_3_88_2/CIN sky130_fd_sc_hd__fa_1
Xrepeater1472 input127/X VGND VGND VPWR VPWR U$$4408/A1 sky130_fd_sc_hd__buf_8
XFILLER_114_944 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1483 U$$3719/A1 VGND VGND VPWR VPWR U$$2623/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_65_0 dadda_fa_5_65_0/A dadda_fa_5_65_0/B dadda_fa_5_65_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_66_0/A dadda_fa_6_65_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1494 U$$4242/B1 VGND VGND VPWR VPWR U$$4516/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_119_1154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_338 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_1108 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_64_8 dadda_fa_1_64_8/A dadda_fa_1_64_8/B dadda_fa_1_64_8/CIN VGND VGND
+ VPWR VPWR dadda_fa_2_65_3/A dadda_fa_3_64_0/A sky130_fd_sc_hd__fa_2
Xdadda_fa_1_57_7 input209/X dadda_fa_1_57_7/B dadda_fa_1_57_7/CIN VGND VGND VPWR VPWR
+ dadda_fa_2_58_2/CIN dadda_fa_2_57_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_279 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_4_0 U$$281/X U$$317/B input201/X VGND VGND VPWR VPWR dadda_fa_7_5_0/B
+ dadda_fa_7_4_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_74_1024 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_196_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_986 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_168_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_210_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_163_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1052 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_90_1 U$$2182/X U$$2315/X U$$2448/X VGND VGND VPWR VPWR dadda_fa_2_91_4/B
+ dadda_fa_2_90_5/B sky130_fd_sc_hd__fa_1
XFILLER_190_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_83_0 U$$1369/Y U$$1503/X U$$1636/X VGND VGND VPWR VPWR dadda_fa_2_84_1/CIN
+ dadda_fa_2_83_4/A sky130_fd_sc_hd__fa_1
XFILLER_116_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4435_1794 VGND VGND VPWR VPWR U$$4435_1794/HI U$$4435/B sky130_fd_sc_hd__conb_1
XFILLER_89_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$4309 U$$4309/A1 U$$4381/A2 U$$4309/B1 U$$4381/B2 VGND VGND VPWR VPWR U$$4310/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3608 input75/X U$$3612/A2 U$$4293/B1 U$$3612/B2 VGND VGND VPWR VPWR U$$3609/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3619 U$$3619/A U$$3623/B VGND VGND VPWR VPWR U$$3619/X sky130_fd_sc_hd__xor2_1
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_35 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2907 U$$30/A1 U$$2995/A2 U$$32/A1 U$$2995/B2 VGND VGND VPWR VPWR U$$2908/A sky130_fd_sc_hd__a22o_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2918 U$$2918/A U$$2920/B VGND VGND VPWR VPWR U$$2918/X sky130_fd_sc_hd__xor2_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _199_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 _209_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XU$$2929 U$$4297/B1 U$$2967/A2 U$$4162/B1 U$$2967/B2 VGND VGND VPWR VPWR U$$2930/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 _215_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 _256_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 _292_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 U$$4011/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 U$$3229/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_364_ _367_/CLK _364_/D VGND VGND VPWR VPWR _364_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_295_ _423_/CLK _295_/D VGND VGND VPWR VPWR _295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_3_114_0_1867 VGND VGND VPWR VPWR dadda_fa_3_114_0/A dadda_fa_3_114_0_1867/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_166_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_6_82_0 dadda_fa_6_82_0/A dadda_fa_6_82_0/B dadda_fa_6_82_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_83_0/B dadda_fa_7_82_0/CIN sky130_fd_sc_hd__fa_1
Xdadda_fa_3_98_0 input254/X dadda_fa_3_98_0/B dadda_fa_3_98_0/CIN VGND VGND VPWR VPWR
+ dadda_fa_4_99_0/B dadda_fa_4_98_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_155_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_190_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_831 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_886 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$380 U$$654/A1 U$$394/A2 U$$654/B1 U$$394/B2 VGND VGND VPWR VPWR U$$381/A sky130_fd_sc_hd__a22o_1
XFILLER_205_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$391 U$$391/A U$$395/B VGND VGND VPWR VPWR U$$391/X sky130_fd_sc_hd__xor2_1
XFILLER_205_583 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_193_939 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_513 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_1033 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_192_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_888 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR _329_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_173_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1280 U$$951/B VGND VGND VPWR VPWR U$$883/B sky130_fd_sc_hd__buf_6
Xrepeater1291 input49/X VGND VGND VPWR VPWR U$$3697/B sky130_fd_sc_hd__buf_8
XFILLER_102_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_925 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_1_62_5 U$$4278/B input215/X dadda_fa_1_62_5/CIN VGND VGND VPWR VPWR dadda_fa_2_63_2/A
+ dadda_fa_2_62_5/A sky130_fd_sc_hd__fa_1
XFILLER_80_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_55_4 U$$2378/X U$$2511/X U$$2644/X VGND VGND VPWR VPWR dadda_fa_2_56_1/CIN
+ dadda_fa_2_55_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_67_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1089 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_48_3 U$$1300/X U$$1433/X U$$1566/X VGND VGND VPWR VPWR dadda_fa_2_49_2/A
+ dadda_fa_2_48_4/CIN sky130_fd_sc_hd__fa_1
XFILLER_82_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_25_2 dadda_fa_4_25_2/A dadda_fa_4_25_2/B dadda_fa_4_25_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_26_0/CIN dadda_fa_5_25_1/CIN sky130_fd_sc_hd__fa_1
Xclkbuf_3_2_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_3_2_0_clk/X sky130_fd_sc_hd__clkbuf_8
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_18_1 input166/X dadda_fa_4_18_1/B dadda_fa_4_18_1/CIN VGND VGND VPWR VPWR
+ dadda_fa_5_19_0/B dadda_fa_5_18_1/B sky130_fd_sc_hd__fa_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$4106 U$$4106/A input55/X VGND VGND VPWR VPWR U$$4106/X sky130_fd_sc_hd__xor2_1
Xdadda_ha_3_21_3 U$$1246/X U$$1379/X VGND VGND VPWR VPWR dadda_fa_4_22_1/B dadda_ha_3_21_3/SUM
+ sky130_fd_sc_hd__ha_1
XFILLER_93_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$4117 U$$4117/A U$$4145/B VGND VGND VPWR VPWR U$$4117/X sky130_fd_sc_hd__xor2_1
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4128 U$$4402/A1 U$$4176/A2 U$$4402/B1 U$$4176/B2 VGND VGND VPWR VPWR U$$4129/A
+ sky130_fd_sc_hd__a22o_1
XU$$4139 U$$4139/A U$$4165/B VGND VGND VPWR VPWR U$$4139/X sky130_fd_sc_hd__xor2_1
XU$$3405 U$$3405/A U$$3424/A VGND VGND VPWR VPWR U$$3405/X sky130_fd_sc_hd__xor2_1
XU$$3416 U$$3416/A1 U$$3416/A2 input122/X U$$3416/B2 VGND VGND VPWR VPWR U$$3417/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_150_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_747 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3427 U$$3510/B VGND VGND VPWR VPWR U$$3427/Y sky130_fd_sc_hd__inv_1
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$3438 U$$3438/A U$$3528/B VGND VGND VPWR VPWR U$$3438/X sky130_fd_sc_hd__xor2_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2704 U$$2704/A U$$2710/B VGND VGND VPWR VPWR U$$2704/X sky130_fd_sc_hd__xor2_1
XU$$3449 U$$3584/B1 U$$3453/A2 U$$3451/A1 U$$3453/B2 VGND VGND VPWR VPWR U$$3450/A
+ sky130_fd_sc_hd__a22o_1
XU$$2715 U$$2715/A1 U$$2737/A2 U$$2717/A1 U$$2737/B2 VGND VGND VPWR VPWR U$$2716/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2726 U$$2726/A U$$2736/B VGND VGND VPWR VPWR U$$2726/X sky130_fd_sc_hd__xor2_1
XFILLER_37_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2737 U$$3557/B1 U$$2737/A2 U$$2737/B1 U$$2737/B2 VGND VGND VPWR VPWR U$$2738/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_20_1 U$$446/X U$$579/X U$$712/X VGND VGND VPWR VPWR dadda_fa_4_21_0/CIN
+ dadda_fa_4_20_2/A sky130_fd_sc_hd__fa_1
XU$$2748 U$$3159/A1 U$$2796/A2 U$$3159/B1 U$$2796/B2 VGND VGND VPWR VPWR U$$2749/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$2759 U$$2759/A U$$2797/B VGND VGND VPWR VPWR U$$2759/X sky130_fd_sc_hd__xor2_1
XFILLER_61_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_416_ _417_/CLK _416_/D VGND VGND VPWR VPWR _416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_347_ _351_/CLK _347_/D VGND VGND VPWR VPWR _347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_278_ _407_/CLK _278_/D VGND VGND VPWR VPWR _278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_72_4 dadda_fa_2_72_4/A dadda_fa_2_72_4/B dadda_fa_2_72_4/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_73_1/CIN dadda_fa_3_72_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_29_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1053 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_636 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_1195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_65_3 dadda_fa_2_65_3/A dadda_fa_2_65_3/B dadda_fa_2_65_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_66_1/B dadda_fa_3_65_3/B sky130_fd_sc_hd__fa_1
Xrepeater903 U$$3922/B1 VGND VGND VPWR VPWR U$$910/A1 sky130_fd_sc_hd__buf_4
XFILLER_151_1048 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater914 U$$2343/A1 VGND VGND VPWR VPWR U$$3028/A1 sky130_fd_sc_hd__clkbuf_4
Xrepeater925 U$$4468/B1 VGND VGND VPWR VPWR U$$3511/A1 sky130_fd_sc_hd__buf_6
Xrepeater936 U$$4055/A1 VGND VGND VPWR VPWR U$$2683/B1 sky130_fd_sc_hd__buf_4
Xdadda_fa_2_58_2 dadda_fa_2_58_2/A dadda_fa_2_58_2/B dadda_fa_2_58_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_59_1/A dadda_fa_3_58_3/A sky130_fd_sc_hd__fa_1
XFILLER_37_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater947 U$$2957/A1 VGND VGND VPWR VPWR U$$4188/B1 sky130_fd_sc_hd__buf_6
XFILLER_65_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater958 input93/X VGND VGND VPWR VPWR U$$4049/B1 sky130_fd_sc_hd__buf_6
XFILLER_37_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrepeater969 U$$4458/A1 VGND VGND VPWR VPWR U$$2951/A1 sky130_fd_sc_hd__buf_4
Xdadda_fa_5_35_1 dadda_fa_5_35_1/A dadda_fa_5_35_1/B dadda_fa_5_35_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_36_0/B dadda_fa_7_35_0/A sky130_fd_sc_hd__fa_1
XFILLER_204_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_28_0 dadda_fa_5_28_0/A dadda_fa_5_28_0/B dadda_fa_5_28_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_29_0/A dadda_fa_6_28_0/CIN sky130_fd_sc_hd__fa_1
XU$$3950 input113/X U$$3968/A2 input114/X U$$3968/B2 VGND VGND VPWR VPWR U$$3951/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$3961 U$$3961/A U$$3967/B VGND VGND VPWR VPWR U$$3961/X sky130_fd_sc_hd__xor2_1
XFILLER_65_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3972 U$$3972/A VGND VGND VPWR VPWR U$$3972/Y sky130_fd_sc_hd__inv_1
XU$$3983 U$$4394/A1 U$$4043/A2 U$$4396/A1 U$$4043/B2 VGND VGND VPWR VPWR U$$3984/A
+ sky130_fd_sc_hd__a22o_1
XU$$3994 U$$3994/A U$$4012/B VGND VGND VPWR VPWR U$$3994/X sky130_fd_sc_hd__xor2_1
XFILLER_91_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$819_1842 VGND VGND VPWR VPWR U$$819_1842/HI U$$819/B1 sky130_fd_sc_hd__conb_1
XFILLER_203_1152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_181_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_102_0 dadda_fa_5_102_0/A dadda_fa_5_102_0/B dadda_fa_5_102_0/CIN VGND
+ VGND VPWR VPWR dadda_fa_6_103_0/A dadda_fa_6_102_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput263 output263/A VGND VGND VPWR VPWR o[105] sky130_fd_sc_hd__buf_2
Xoutput274 output274/A VGND VGND VPWR VPWR o[115] sky130_fd_sc_hd__buf_2
XFILLER_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput285 output285/A VGND VGND VPWR VPWR o[125] sky130_fd_sc_hd__buf_2
XFILLER_173_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput296 output296/A VGND VGND VPWR VPWR o[1] sky130_fd_sc_hd__buf_2
XFILLER_59_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_1178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_199_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_1_60_2 U$$2787/X U$$2920/X U$$3053/X VGND VGND VPWR VPWR dadda_fa_2_61_1/A
+ dadda_fa_2_60_4/A sky130_fd_sc_hd__fa_1
XFILLER_102_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_639 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_53_1 U$$778/X U$$911/X U$$1044/X VGND VGND VPWR VPWR dadda_fa_2_54_0/CIN
+ dadda_fa_2_53_3/CIN sky130_fd_sc_hd__fa_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_4_30_0 dadda_fa_4_30_0/A dadda_fa_4_30_0/B dadda_fa_4_30_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_31_0/A dadda_fa_5_30_1/A sky130_fd_sc_hd__fa_1
XFILLER_56_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_1_46_0 U$$99/X U$$232/X U$$365/X VGND VGND VPWR VPWR dadda_fa_2_47_1/CIN
+ dadda_fa_2_46_4/A sky130_fd_sc_hd__fa_1
XFILLER_71_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_203_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_1244 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_201_ _329_/CLK _201_/D VGND VGND VPWR VPWR _201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_211_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$1104 final_adder.U$$174/A final_adder.U$$883/X VGND VGND VPWR VPWR
+ output363/A sky130_fd_sc_hd__xor2_1
XFILLER_168_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_949 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1115 final_adder.U$$164/B final_adder.U$$935/X VGND VGND VPWR VPWR
+ output375/A sky130_fd_sc_hd__xor2_1
XFILLER_17_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1126 final_adder.U$$152/A final_adder.U$$861/X VGND VGND VPWR VPWR
+ output260/A sky130_fd_sc_hd__xor2_2
XFILLER_99_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$1137 final_adder.U$$142/B final_adder.U$$913/X VGND VGND VPWR VPWR
+ output272/A sky130_fd_sc_hd__xor2_1
XFILLER_104_1061 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$1148 final_adder.U$$130/A final_adder.U$$839/X VGND VGND VPWR VPWR
+ output284/A sky130_fd_sc_hd__xor2_1
XFILLER_99_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_3_82_3 dadda_fa_3_82_3/A dadda_fa_3_82_3/B dadda_fa_3_82_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_83_1/B dadda_fa_4_82_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_178_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_75_2 dadda_fa_3_75_2/A dadda_fa_3_75_2/B dadda_fa_3_75_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_76_1/A dadda_fa_4_75_2/B sky130_fd_sc_hd__fa_1
XFILLER_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_68_1 dadda_fa_3_68_1/A dadda_fa_3_68_1/B dadda_fa_3_68_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_69_0/CIN dadda_fa_4_68_2/A sky130_fd_sc_hd__fa_1
XFILLER_78_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_6_45_0 dadda_fa_6_45_0/A dadda_fa_6_45_0/B dadda_fa_6_45_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_7_46_0/B dadda_fa_7_45_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_78_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$3202 U$$3202/A U$$3208/B VGND VGND VPWR VPWR U$$3202/X sky130_fd_sc_hd__xor2_1
XFILLER_171_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3213 U$$610/A1 U$$3229/A2 U$$3213/B1 U$$3227/B2 VGND VGND VPWR VPWR U$$3214/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3224 U$$3224/A U$$3288/A VGND VGND VPWR VPWR U$$3224/X sky130_fd_sc_hd__xor2_1
XU$$3235 U$$3235/A1 U$$3241/A2 U$$3235/B1 U$$3241/B2 VGND VGND VPWR VPWR U$$3236/A
+ sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$17 _313_/Q _185_/Q VGND VGND VPWR VPWR final_adder.U$$239/B1 final_adder.U$$238/B
+ sky130_fd_sc_hd__ha_1
XU$$2501 U$$2501/A U$$2597/B VGND VGND VPWR VPWR U$$2501/X sky130_fd_sc_hd__xor2_1
XFILLER_46_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$28 _324_/Q _196_/Q VGND VGND VPWR VPWR final_adder.U$$997/B1 final_adder.U$$226/A
+ sky130_fd_sc_hd__ha_1
XU$$3246 U$$3246/A U$$3288/A VGND VGND VPWR VPWR U$$3246/X sky130_fd_sc_hd__xor2_1
XFILLER_111_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3257 U$$517/A1 U$$3263/A2 U$$517/B1 U$$3263/B2 VGND VGND VPWR VPWR U$$3258/A sky130_fd_sc_hd__a22o_1
XU$$2512 U$$44/B1 U$$2596/A2 U$$3882/B1 U$$2596/B2 VGND VGND VPWR VPWR U$$2513/A sky130_fd_sc_hd__a22o_1
Xdadda_fa_4_104_2 dadda_fa_4_104_2/A dadda_fa_4_104_2/B dadda_fa_4_104_2/CIN VGND
+ VGND VPWR VPWR dadda_fa_5_105_0/CIN dadda_fa_5_104_1/CIN sky130_fd_sc_hd__fa_1
XU$$3268 U$$3268/A U$$3286/B VGND VGND VPWR VPWR U$$3268/X sky130_fd_sc_hd__xor2_1
Xfinal_adder.U$$39 _335_/Q _207_/Q VGND VGND VPWR VPWR final_adder.U$$217/B1 final_adder.U$$216/B
+ sky130_fd_sc_hd__ha_1
XU$$2523 U$$2523/A U$$2543/B VGND VGND VPWR VPWR U$$2523/X sky130_fd_sc_hd__xor2_1
XU$$3279 U$$3414/B1 U$$3285/A2 U$$3281/A1 U$$3285/B2 VGND VGND VPWR VPWR U$$3280/A
+ sky130_fd_sc_hd__a22o_1
XU$$2534 U$$3902/B1 U$$2576/A2 U$$2808/B1 U$$2576/B2 VGND VGND VPWR VPWR U$$2535/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2545 U$$2545/A U$$2569/B VGND VGND VPWR VPWR U$$2545/X sky130_fd_sc_hd__xor2_1
XU$$1800 U$$1800/A U$$1832/B VGND VGND VPWR VPWR U$$1800/X sky130_fd_sc_hd__xor2_1
XU$$2556 U$$4335/B1 U$$2588/A2 U$$366/A1 U$$2588/B2 VGND VGND VPWR VPWR U$$2557/A
+ sky130_fd_sc_hd__a22o_1
XU$$1811 U$$989/A1 U$$1831/A2 U$$991/A1 U$$1831/B2 VGND VGND VPWR VPWR U$$1812/A sky130_fd_sc_hd__a22o_1
XFILLER_94_1049 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_206_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1822 U$$1822/A U$$1870/B VGND VGND VPWR VPWR U$$1822/X sky130_fd_sc_hd__xor2_1
XFILLER_61_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$2567 U$$2567/A U$$2569/B VGND VGND VPWR VPWR U$$2567/X sky130_fd_sc_hd__xor2_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$2578 U$$934/A1 U$$2470/X U$$936/A1 U$$2471/X VGND VGND VPWR VPWR U$$2579/A sky130_fd_sc_hd__a22o_1
XU$$1833 U$$52/A1 U$$1839/A2 U$$52/B1 U$$1839/B2 VGND VGND VPWR VPWR U$$1834/A sky130_fd_sc_hd__a22o_1
XU$$2589 U$$2589/A U$$2602/A VGND VGND VPWR VPWR U$$2589/X sky130_fd_sc_hd__xor2_1
XU$$1844 U$$1844/A U$$1880/B VGND VGND VPWR VPWR U$$1844/X sky130_fd_sc_hd__xor2_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1855 U$$483/B1 U$$1879/A2 U$$76/A1 U$$1879/B2 VGND VGND VPWR VPWR U$$1856/A sky130_fd_sc_hd__a22o_1
XU$$1866 U$$1866/A U$$1912/B VGND VGND VPWR VPWR U$$1866/X sky130_fd_sc_hd__xor2_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1877 U$$2425/A1 U$$1877/A2 U$$2016/A1 U$$1877/B2 VGND VGND VPWR VPWR U$$1878/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_271 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1888 U$$1888/A U$$1917/A VGND VGND VPWR VPWR U$$1888/X sky130_fd_sc_hd__xor2_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$1899 U$$2445/B1 U$$1913/A2 U$$2312/A1 U$$1903/B2 VGND VGND VPWR VPWR U$$1900/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_7_118_0 dadda_fa_7_118_0/A dadda_fa_7_118_0/B dadda_fa_7_118_0/CIN VGND
+ VGND VPWR VPWR _415_/D _286_/D sky130_fd_sc_hd__fa_1
XFILLER_147_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_183_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_644 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_157_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_70_1 dadda_fa_2_70_1/A dadda_fa_2_70_1/B dadda_fa_2_70_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_71_0/CIN dadda_fa_3_70_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_69_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdadda_fa_2_63_0 dadda_fa_2_63_0/A dadda_fa_2_63_0/B dadda_fa_2_63_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_64_0/B dadda_fa_3_63_2/B sky130_fd_sc_hd__fa_1
XFILLER_111_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater700 U$$3978/X VGND VGND VPWR VPWR U$$4101/B2 sky130_fd_sc_hd__buf_6
Xrepeater711 U$$3777/B2 VGND VGND VPWR VPWR U$$3753/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$518 final_adder.U$$526/B final_adder.U$$518/B VGND VGND VPWR VPWR
+ final_adder.U$$638/B sky130_fd_sc_hd__and2_1
Xrepeater722 U$$3696/B2 VGND VGND VPWR VPWR U$$3686/B2 sky130_fd_sc_hd__buf_6
Xfinal_adder.U$$529 final_adder.U$$528/B final_adder.U$$413/X final_adder.U$$405/X
+ VGND VGND VPWR VPWR final_adder.U$$529/X sky130_fd_sc_hd__a21o_1
XFILLER_42_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater733 U$$3430/X VGND VGND VPWR VPWR U$$3517/B2 sky130_fd_sc_hd__buf_6
XFILLER_85_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater744 U$$3156/X VGND VGND VPWR VPWR U$$3241/B2 sky130_fd_sc_hd__buf_6
XFILLER_96_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater755 U$$3118/B2 VGND VGND VPWR VPWR U$$3132/B2 sky130_fd_sc_hd__buf_4
Xrepeater766 U$$396/B2 VGND VGND VPWR VPWR U$$350/B2 sky130_fd_sc_hd__buf_6
Xrepeater777 U$$2828/B2 VGND VGND VPWR VPWR U$$2782/B2 sky130_fd_sc_hd__buf_4
XU$$4470 input97/X U$$4388/X input99/X U$$4486/B2 VGND VGND VPWR VPWR U$$4471/A sky130_fd_sc_hd__a22o_1
Xrepeater788 U$$2737/B2 VGND VGND VPWR VPWR U$$2735/B2 sky130_fd_sc_hd__buf_4
Xrepeater799 U$$2403/B2 VGND VGND VPWR VPWR U$$2359/B2 sky130_fd_sc_hd__clkbuf_4
XU$$4481 U$$4481/A U$$4481/B VGND VGND VPWR VPWR U$$4481/X sky130_fd_sc_hd__xor2_1
XU$$4492 U$$4492/A1 U$$4388/X U$$4494/A1 U$$4494/B2 VGND VGND VPWR VPWR U$$4493/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$3780 U$$3780/A U$$3834/B VGND VGND VPWR VPWR U$$3780/X sky130_fd_sc_hd__xor2_1
XFILLER_44_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3791 U$$4476/A1 U$$3793/A2 U$$4476/B1 U$$3793/B2 VGND VGND VPWR VPWR U$$3792/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_178_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_1037 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_165_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdadda_fa_4_92_2 dadda_fa_4_92_2/A dadda_fa_4_92_2/B dadda_fa_4_92_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_93_0/CIN dadda_fa_5_92_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_4_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_22 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_4_85_1 dadda_fa_4_85_1/A dadda_fa_4_85_1/B dadda_fa_4_85_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_86_0/B dadda_fa_5_85_1/B sky130_fd_sc_hd__fa_1
XFILLER_118_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_7_62_0 dadda_fa_7_62_0/A dadda_fa_7_62_0/B dadda_fa_7_62_0/CIN VGND VGND
+ VPWR VPWR _359_/D _230_/D sky130_fd_sc_hd__fa_1
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_4_78_0 dadda_fa_4_78_0/A dadda_fa_4_78_0/B dadda_fa_4_78_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_79_0/A dadda_fa_5_78_1/A sky130_fd_sc_hd__fa_1
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_937 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$902 U$$902/A1 U$$906/A2 U$$82/A1 U$$906/B2 VGND VGND VPWR VPWR U$$903/A sky130_fd_sc_hd__a22o_1
XU$$913 U$$913/A U$$919/B VGND VGND VPWR VPWR U$$913/X sky130_fd_sc_hd__xor2_1
XFILLER_21_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$924 U$$924/A1 U$$950/A2 U$$926/A1 U$$950/B2 VGND VGND VPWR VPWR U$$925/A sky130_fd_sc_hd__a22o_1
XFILLER_84_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$935 U$$935/A U$$959/A VGND VGND VPWR VPWR U$$935/X sky130_fd_sc_hd__xor2_1
XFILLER_62_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XU$$946 U$$946/A1 U$$826/X U$$948/A1 U$$827/X VGND VGND VPWR VPWR U$$947/A sky130_fd_sc_hd__a22o_1
XFILLER_204_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$957 U$$957/A U$$958/A VGND VGND VPWR VPWR U$$957/X sky130_fd_sc_hd__xor2_1
XFILLER_189_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$968 U$$968/A U$$968/B VGND VGND VPWR VPWR U$$968/X sky130_fd_sc_hd__xor2_1
XU$$1107 U$$1107/A U$$1139/B VGND VGND VPWR VPWR U$$1107/X sky130_fd_sc_hd__xor2_1
XFILLER_16_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$979 U$$979/A1 U$$979/A2 U$$22/A1 U$$979/B2 VGND VGND VPWR VPWR U$$980/A sky130_fd_sc_hd__a22o_1
XU$$1118 U$$1666/A1 U$$1136/A2 U$$1666/B1 U$$1136/B2 VGND VGND VPWR VPWR U$$1119/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1129 U$$1129/A U$$1137/B VGND VGND VPWR VPWR U$$1129/X sky130_fd_sc_hd__xor2_1
XFILLER_203_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_203_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_1093 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_961 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_172_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_184_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_953 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_3_80_0 dadda_fa_3_80_0/A dadda_fa_3_80_0/B dadda_fa_3_80_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_81_0/B dadda_fa_4_80_1/CIN sky130_fd_sc_hd__fa_1
XFILLER_124_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_915 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_872 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_208_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$3010 U$$3010/A U$$3013/A VGND VGND VPWR VPWR U$$3010/X sky130_fd_sc_hd__xor2_1
Xdadda_fa_2_42_5 dadda_fa_2_42_5/A dadda_fa_2_42_5/B dadda_fa_2_42_5/CIN VGND VGND
+ VPWR VPWR dadda_fa_3_43_2/A dadda_fa_4_42_0/A sky130_fd_sc_hd__fa_1
XU$$3021 U$$3021/A U$$3075/B VGND VGND VPWR VPWR U$$3021/X sky130_fd_sc_hd__xor2_1
XU$$3032 U$$3032/A1 U$$3082/A2 U$$4404/A1 U$$3082/B2 VGND VGND VPWR VPWR U$$3033/A
+ sky130_fd_sc_hd__a22o_1
XU$$3043 U$$3043/A U$$3125/B VGND VGND VPWR VPWR U$$3043/X sky130_fd_sc_hd__xor2_1
XFILLER_75_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$3054 U$$4424/A1 U$$3060/A2 U$$3876/B1 U$$3060/B2 VGND VGND VPWR VPWR U$$3055/A
+ sky130_fd_sc_hd__a22o_1
XU$$2320 U$$3416/A1 U$$2326/A2 U$$3829/A1 U$$2326/B2 VGND VGND VPWR VPWR U$$2321/A
+ sky130_fd_sc_hd__a22o_1
XU$$3065 U$$3065/A U$$3109/B VGND VGND VPWR VPWR U$$3065/X sky130_fd_sc_hd__xor2_1
XFILLER_62_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_35_4 U$$1939/X U$$2072/X U$$2205/X VGND VGND VPWR VPWR dadda_fa_3_36_1/CIN
+ dadda_fa_3_35_3/CIN sky130_fd_sc_hd__fa_1
XU$$2331 input29/X VGND VGND VPWR VPWR U$$2331/Y sky130_fd_sc_hd__inv_1
XU$$3076 U$$3211/B1 U$$3098/A2 U$$3352/A1 U$$3098/B2 VGND VGND VPWR VPWR U$$3077/A
+ sky130_fd_sc_hd__a22o_1
XU$$3087 U$$3087/A U$$3117/B VGND VGND VPWR VPWR U$$3087/X sky130_fd_sc_hd__xor2_1
XU$$2342 U$$2342/A U$$2366/B VGND VGND VPWR VPWR U$$2342/X sky130_fd_sc_hd__xor2_1
XFILLER_207_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$2353 U$$2625/B1 U$$2359/A2 U$$2492/A1 U$$2359/B2 VGND VGND VPWR VPWR U$$2354/A
+ sky130_fd_sc_hd__a22o_1
XU$$3098 U$$3644/B1 U$$3098/A2 U$$3511/A1 U$$3098/B2 VGND VGND VPWR VPWR U$$3099/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2364 U$$2364/A U$$2366/B VGND VGND VPWR VPWR U$$2364/X sky130_fd_sc_hd__xor2_1
XU$$2375 U$$3880/B1 U$$2463/A2 U$$3882/B1 U$$2463/B2 VGND VGND VPWR VPWR U$$2376/A
+ sky130_fd_sc_hd__a22o_1
XU$$1630 U$$1630/A U$$1638/B VGND VGND VPWR VPWR U$$1630/X sky130_fd_sc_hd__xor2_1
XFILLER_22_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1641 U$$4516/B1 U$$1511/X U$$1641/B1 U$$1512/X VGND VGND VPWR VPWR U$$1642/A sky130_fd_sc_hd__a22o_1
XFILLER_34_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2386 U$$2386/A U$$2426/B VGND VGND VPWR VPWR U$$2386/X sky130_fd_sc_hd__xor2_1
XU$$2397 U$$3902/B1 U$$2403/A2 U$$2808/B1 U$$2403/B2 VGND VGND VPWR VPWR U$$2398/A
+ sky130_fd_sc_hd__a22o_1
XU$$1652 U$$2198/B1 U$$1696/A2 U$$2063/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1653/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$1663 U$$1663/A U$$1679/B VGND VGND VPWR VPWR U$$1663/X sky130_fd_sc_hd__xor2_1
XFILLER_210_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1674 U$$989/A1 U$$1696/A2 U$$991/A1 U$$1696/B2 VGND VGND VPWR VPWR U$$1675/A sky130_fd_sc_hd__a22o_1
XU$$1685 U$$1685/A U$$1689/B VGND VGND VPWR VPWR U$$1685/X sky130_fd_sc_hd__xor2_1
XU$$1696 U$$3612/B1 U$$1696/A2 U$$874/B1 U$$1696/B2 VGND VGND VPWR VPWR U$$1697/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_1106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_95_0 dadda_fa_5_95_0/A dadda_fa_5_95_0/B dadda_fa_5_95_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_96_0/A dadda_fa_6_95_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_162_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$304 final_adder.U$$306/B final_adder.U$$304/B VGND VGND VPWR VPWR
+ final_adder.U$$430/B sky130_fd_sc_hd__and2_1
Xfinal_adder.U$$315 final_adder.U$$314/B final_adder.U$$189/X final_adder.U$$187/X
+ VGND VGND VPWR VPWR final_adder.U$$315/X sky130_fd_sc_hd__a21o_1
Xfinal_adder.U$$326 final_adder.U$$328/B final_adder.U$$326/B VGND VGND VPWR VPWR
+ final_adder.U$$452/B sky130_fd_sc_hd__and2_1
XU$$4_1758 VGND VGND VPWR VPWR U$$4_1758/HI U$$4/A3 sky130_fd_sc_hd__conb_1
XFILLER_85_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater530 U$$2828/A2 VGND VGND VPWR VPWR U$$2782/A2 sky130_fd_sc_hd__buf_4
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfinal_adder.U$$337 final_adder.U$$336/B final_adder.U$$211/X final_adder.U$$209/X
+ VGND VGND VPWR VPWR final_adder.U$$337/X sky130_fd_sc_hd__a21o_1
Xrepeater541 U$$2737/A2 VGND VGND VPWR VPWR U$$2735/A2 sky130_fd_sc_hd__buf_4
XTAP_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$348 final_adder.U$$350/B final_adder.U$$348/B VGND VGND VPWR VPWR
+ final_adder.U$$474/B sky130_fd_sc_hd__and2_1
XTAP_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater552 U$$2403/A2 VGND VGND VPWR VPWR U$$2359/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_84_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfinal_adder.U$$359 final_adder.U$$358/B final_adder.U$$233/X final_adder.U$$231/X
+ VGND VGND VPWR VPWR final_adder.U$$359/X sky130_fd_sc_hd__a21o_1
Xrepeater563 U$$2326/A2 VGND VGND VPWR VPWR U$$2284/A2 sky130_fd_sc_hd__buf_4
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater574 U$$2059/X VGND VGND VPWR VPWR U$$2169/A2 sky130_fd_sc_hd__buf_6
XU$$209 U$$72/A1 U$$209/A2 U$$74/A1 U$$209/B2 VGND VGND VPWR VPWR U$$210/A sky130_fd_sc_hd__a22o_1
XFILLER_211_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater585 U$$1785/X VGND VGND VPWR VPWR U$$1869/A2 sky130_fd_sc_hd__clkbuf_8
Xrepeater596 U$$1746/A2 VGND VGND VPWR VPWR U$$1750/A2 sky130_fd_sc_hd__buf_4
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_197_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_1009 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_200_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_205_1077 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_194_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1109 input75/X VGND VGND VPWR VPWR U$$4430/A1 sky130_fd_sc_hd__buf_6
XFILLER_107_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_111_2 U$$4086/X U$$4219/X U$$4352/X VGND VGND VPWR VPWR dadda_fa_4_112_1/CIN
+ dadda_fa_4_111_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_135_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_3_104_1 U$$4205/X U$$4338/X U$$4471/X VGND VGND VPWR VPWR dadda_fa_4_105_0/CIN
+ dadda_fa_4_104_2/A sky130_fd_sc_hd__fa_1
XFILLER_162_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_986 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_699 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_1149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_6_125_0 input157/X dadda_fa_6_125_0/B dadda_fa_6_125_0/CIN VGND VGND VPWR
+ VPWR dadda_fa_7_126_0/B dadda_fa_7_125_0/CIN sky130_fd_sc_hd__fa_1
XTAP_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_0_68_4 U$$1872/X U$$2005/X U$$2138/X VGND VGND VPWR VPWR dadda_fa_1_69_7/A
+ dadda_fa_1_68_8/CIN sky130_fd_sc_hd__fa_1
XFILLER_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_45_3 dadda_fa_3_45_3/A dadda_fa_3_45_3/B dadda_fa_3_45_3/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_46_1/B dadda_fa_4_45_2/CIN sky130_fd_sc_hd__fa_1
XTAP_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$871 final_adder.U$$774/X final_adder.U$$727/X final_adder.U$$775/X
+ VGND VGND VPWR VPWR final_adder.U$$871/X sky130_fd_sc_hd__a21o_1
XU$$710 U$$710/A U$$712/B VGND VGND VPWR VPWR U$$710/X sky130_fd_sc_hd__xor2_1
XFILLER_17_812 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_38_2 dadda_fa_3_38_2/A dadda_fa_3_38_2/B dadda_fa_3_38_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_39_1/A dadda_fa_4_38_2/B sky130_fd_sc_hd__fa_1
XFILLER_91_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$721 U$$995/A1 U$$739/A2 U$$721/B1 U$$739/B2 VGND VGND VPWR VPWR U$$722/A sky130_fd_sc_hd__a22o_1
Xfinal_adder.U$$893 final_adder.U$$796/X final_adder.U$$505/X final_adder.U$$797/X
+ VGND VGND VPWR VPWR final_adder.U$$893/X sky130_fd_sc_hd__a21o_1
XFILLER_28_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$732 U$$732/A U$$740/B VGND VGND VPWR VPWR U$$732/X sky130_fd_sc_hd__xor2_1
XFILLER_112_1182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$743 U$$878/B1 U$$749/A2 U$$745/A1 U$$749/B2 VGND VGND VPWR VPWR U$$744/A sky130_fd_sc_hd__a22o_1
XU$$754 U$$754/A U$$796/B VGND VGND VPWR VPWR U$$754/X sky130_fd_sc_hd__xor2_1
XFILLER_186_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$765 U$$80/A1 U$$793/A2 U$$82/A1 U$$793/B2 VGND VGND VPWR VPWR U$$766/A sky130_fd_sc_hd__a22o_1
XU$$776 U$$776/A U$$784/B VGND VGND VPWR VPWR U$$776/X sky130_fd_sc_hd__xor2_1
XFILLER_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$787 U$$787/A1 U$$793/A2 U$$926/A1 U$$793/B2 VGND VGND VPWR VPWR U$$788/A sky130_fd_sc_hd__a22o_1
XU$$798 U$$798/A U$$808/B VGND VGND VPWR VPWR U$$798/X sky130_fd_sc_hd__xor2_1
XFILLER_31_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_1161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1610 input111/X VGND VGND VPWR VPWR U$$4494/A1 sky130_fd_sc_hd__buf_4
XANTENNA_4 _327_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater1621 U$$1330/B VGND VGND VPWR VPWR U$$1286/B sky130_fd_sc_hd__buf_6
Xrepeater1632 input109/X VGND VGND VPWR VPWR U$$3578/A1 sky130_fd_sc_hd__buf_4
Xrepeater1643 U$$4490/A1 VGND VGND VPWR VPWR U$$517/A1 sky130_fd_sc_hd__buf_6
XFILLER_141_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater1654 U$$650/A1 VGND VGND VPWR VPWR U$$787/A1 sky130_fd_sc_hd__buf_8
Xrepeater1665 U$$2701/B1 VGND VGND VPWR VPWR U$$2975/B1 sky130_fd_sc_hd__buf_6
Xrepeater1676 input104/X VGND VGND VPWR VPWR U$$4480/B1 sky130_fd_sc_hd__buf_6
XFILLER_154_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater1687 U$$4478/A1 VGND VGND VPWR VPWR U$$4476/B1 sky130_fd_sc_hd__buf_6
Xrepeater1698 U$$3517/A1 VGND VGND VPWR VPWR U$$3243/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_101_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_ha_2_27_2 U$$859/X U$$992/X VGND VGND VPWR VPWR dadda_fa_3_28_2/CIN dadda_fa_4_27_0/A
+ sky130_fd_sc_hd__ha_1
XFILLER_94_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdadda_fa_2_40_2 U$$2348/X U$$2481/X U$$2614/X VGND VGND VPWR VPWR dadda_fa_3_41_1/A
+ dadda_fa_3_40_3/A sky130_fd_sc_hd__fa_1
XFILLER_48_981 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_1047 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_940 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_207_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_2_33_1 U$$472/X U$$605/X U$$738/X VGND VGND VPWR VPWR dadda_fa_3_34_0/CIN
+ dadda_fa_3_33_2/CIN sky130_fd_sc_hd__fa_1
XFILLER_19_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_962 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_179_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_5_10_0 U$$692/X U$$712/B input140/X VGND VGND VPWR VPWR dadda_fa_6_11_0/A
+ dadda_fa_6_10_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2150 U$$2150/A U$$2150/B VGND VGND VPWR VPWR U$$2150/X sky130_fd_sc_hd__xor2_1
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_26_0 U$$59/X U$$192/X U$$325/X VGND VGND VPWR VPWR dadda_fa_3_27_2/B dadda_fa_3_26_3/B
+ sky130_fd_sc_hd__fa_2
XFILLER_63_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XU$$2161 U$$2981/B1 U$$2183/A2 U$$2848/A1 U$$2183/B2 VGND VGND VPWR VPWR U$$2162/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$2172 U$$2172/A U$$2178/B VGND VGND VPWR VPWR U$$2172/X sky130_fd_sc_hd__xor2_1
XFILLER_35_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$2183 U$$4099/B1 U$$2183/A2 U$$4375/B1 U$$2183/B2 VGND VGND VPWR VPWR U$$2184/A
+ sky130_fd_sc_hd__a22o_1
XU$$2194 U$$2311/B VGND VGND VPWR VPWR U$$2194/Y sky130_fd_sc_hd__inv_1
XFILLER_23_859 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$1460 U$$90/A1 U$$1470/A2 U$$92/A1 U$$1470/B2 VGND VGND VPWR VPWR U$$1461/A sky130_fd_sc_hd__a22o_1
XFILLER_50_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_195_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XU$$1471 U$$1471/A U$$1506/A VGND VGND VPWR VPWR U$$1471/X sky130_fd_sc_hd__xor2_1
XFILLER_37_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XU$$1482 U$$660/A1 U$$1504/A2 U$$2717/A1 U$$1504/B2 VGND VGND VPWR VPWR U$$1483/A
+ sky130_fd_sc_hd__a22o_1
XU$$1493 U$$1493/A U$$1499/B VGND VGND VPWR VPWR U$$1493/X sky130_fd_sc_hd__xor2_1
XFILLER_194_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_1121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_175_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1201 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_191_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_945 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_85_4 U$$3103/X U$$3236/X U$$3369/X VGND VGND VPWR VPWR dadda_fa_2_86_3/CIN
+ dadda_fa_2_85_5/CIN sky130_fd_sc_hd__fa_1
XFILLER_103_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_1_78_3 U$$2424/X U$$2557/X U$$2690/X VGND VGND VPWR VPWR dadda_fa_2_79_1/B
+ dadda_fa_2_78_4/B sky130_fd_sc_hd__fa_1
XFILLER_44_1010 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_4_55_2 dadda_fa_4_55_2/A dadda_fa_4_55_2/B dadda_fa_4_55_2/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_56_0/CIN dadda_fa_5_55_1/CIN sky130_fd_sc_hd__fa_1
XTAP_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$101 _397_/Q _269_/Q VGND VGND VPWR VPWR final_adder.U$$155/B1 final_adder.U$$154/B
+ sky130_fd_sc_hd__ha_1
XTAP_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$112 _408_/Q _280_/Q VGND VGND VPWR VPWR final_adder.U$$913/B1 final_adder.U$$142/A
+ sky130_fd_sc_hd__ha_1
XTAP_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$123 _419_/Q _291_/Q VGND VGND VPWR VPWR final_adder.U$$133/B1 final_adder.U$$132/B
+ sky130_fd_sc_hd__ha_1
XTAP_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_4_48_1 dadda_fa_4_48_1/A dadda_fa_4_48_1/B dadda_fa_4_48_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_5_49_0/B dadda_fa_5_48_1/B sky130_fd_sc_hd__fa_1
XFILLER_66_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfinal_adder.U$$134 final_adder.U$$134/A final_adder.U$$134/B VGND VGND VPWR VPWR
+ final_adder.U$$262/B sky130_fd_sc_hd__and2_1
XTAP_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$145 final_adder.U$$144/B final_adder.U$$915/B1 final_adder.U$$145/B1
+ VGND VGND VPWR VPWR final_adder.U$$145/X sky130_fd_sc_hd__a21o_1
XTAP_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_7_25_0 dadda_fa_7_25_0/A dadda_fa_7_25_0/B dadda_fa_7_25_0/CIN VGND VGND
+ VPWR VPWR _322_/D _193_/D sky130_fd_sc_hd__fa_2
Xfinal_adder.U$$156 final_adder.U$$156/A final_adder.U$$156/B VGND VGND VPWR VPWR
+ final_adder.U$$284/B sky130_fd_sc_hd__and2_1
XTAP_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfinal_adder.U$$167 final_adder.U$$166/B final_adder.U$$937/B1 final_adder.U$$167/B1
+ VGND VGND VPWR VPWR final_adder.U$$167/X sky130_fd_sc_hd__a21o_1
XTAP_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfinal_adder.U$$178 final_adder.U$$178/A final_adder.U$$178/B VGND VGND VPWR VPWR
+ final_adder.U$$306/B sky130_fd_sc_hd__and2_1
XTAP_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$189 final_adder.U$$188/B final_adder.U$$959/B1 final_adder.U$$189/B1
+ VGND VGND VPWR VPWR final_adder.U$$189/X sky130_fd_sc_hd__a21o_1
Xrepeater393 U$$882/A2 VGND VGND VPWR VPWR U$$872/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_202_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_198_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_380_ _380_/CLK _380_/D VGND VGND VPWR VPWR _380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_892 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_167_864 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_0_73_2 U$$1483/X U$$1616/X U$$1749/X VGND VGND VPWR VPWR dadda_fa_1_74_8/A
+ dadda_fa_2_73_0/A sky130_fd_sc_hd__fa_1
XFILLER_27_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput130 c[100] VGND VGND VPWR VPWR input130/X sky130_fd_sc_hd__buf_4
XFILLER_49_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput141 c[110] VGND VGND VPWR VPWR input141/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_3_50_1 dadda_fa_3_50_1/A dadda_fa_3_50_1/B dadda_fa_3_50_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_51_0/CIN dadda_fa_4_50_2/A sky130_fd_sc_hd__fa_1
Xinput152 c[120] VGND VGND VPWR VPWR input152/X sky130_fd_sc_hd__clkbuf_4
Xdadda_fa_0_66_1 U$$538/X U$$671/X U$$804/X VGND VGND VPWR VPWR dadda_fa_1_67_5/CIN
+ dadda_fa_1_66_7/CIN sky130_fd_sc_hd__fa_1
Xinput163 c[15] VGND VGND VPWR VPWR input163/X sky130_fd_sc_hd__clkbuf_4
XTAP_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdadda_fa_3_43_0 dadda_fa_3_43_0/A dadda_fa_3_43_0/B dadda_fa_3_43_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_4_44_0/B dadda_fa_4_43_1/CIN sky130_fd_sc_hd__fa_1
Xinput174 c[25] VGND VGND VPWR VPWR input174/X sky130_fd_sc_hd__clkbuf_2
Xinput185 c[35] VGND VGND VPWR VPWR input185/X sky130_fd_sc_hd__buf_2
XTAP_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput196 c[45] VGND VGND VPWR VPWR input196/X sky130_fd_sc_hd__clkbuf_1
Xdadda_fa_0_59_0 U$$125/X U$$258/X U$$391/X VGND VGND VPWR VPWR dadda_fa_1_60_6/B
+ dadda_fa_1_59_8/A sky130_fd_sc_hd__fa_1
XFILLER_97_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfinal_adder.U$$690 final_adder.U$$706/B final_adder.U$$690/B VGND VGND VPWR VPWR
+ final_adder.U$$770/A sky130_fd_sc_hd__and2_1
XTAP_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$540 U$$540/A U$$546/B VGND VGND VPWR VPWR U$$540/X sky130_fd_sc_hd__xor2_1
XTAP_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XU$$551 U$$685/A U$$551/B VGND VGND VPWR VPWR U$$551/X sky130_fd_sc_hd__and2_1
XU$$562 U$$836/A1 U$$578/A2 U$$975/A1 U$$578/B2 VGND VGND VPWR VPWR U$$563/A sky130_fd_sc_hd__a22o_1
XTAP_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$573 U$$573/A U$$607/B VGND VGND VPWR VPWR U$$573/X sky130_fd_sc_hd__xor2_1
XU$$584 U$$36/A1 U$$606/A2 U$$38/A1 U$$606/B2 VGND VGND VPWR VPWR U$$585/A sky130_fd_sc_hd__a22o_1
XFILLER_205_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_189_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_204_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XU$$595 U$$595/A U$$625/B VGND VGND VPWR VPWR U$$595/X sky130_fd_sc_hd__xor2_1
XFILLER_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XU$$956_1844 VGND VGND VPWR VPWR U$$956_1844/HI U$$956/B1 sky130_fd_sc_hd__conb_1
XFILLER_32_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_7_100_0 dadda_fa_7_100_0/A dadda_fa_7_100_0/B dadda_fa_7_100_0/CIN VGND
+ VGND VPWR VPWR _397_/D _268_/D sky130_fd_sc_hd__fa_1
XFILLER_173_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XU$$4493_1823 VGND VGND VPWR VPWR U$$4493_1823/HI U$$4493/B sky130_fd_sc_hd__conb_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_173_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdadda_fa_2_95_3 U$$3788/X U$$3921/X U$$4054/X VGND VGND VPWR VPWR dadda_fa_3_96_1/B
+ dadda_fa_3_95_3/B sky130_fd_sc_hd__fa_1
XFILLER_172_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1440 U$$1638/B VGND VGND VPWR VPWR U$$1628/B sky130_fd_sc_hd__buf_6
XFILLER_99_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrepeater1451 U$$1449/B VGND VGND VPWR VPWR U$$1405/B sky130_fd_sc_hd__buf_6
XFILLER_67_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdadda_fa_2_88_2 U$$4306/X U$$4439/X input243/X VGND VGND VPWR VPWR dadda_fa_3_89_1/A
+ dadda_fa_3_88_3/A sky130_fd_sc_hd__fa_1
Xrepeater1462 U$$4408/B1 VGND VGND VPWR VPWR U$$4273/A1 sky130_fd_sc_hd__buf_6
XFILLER_113_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1473 U$$3447/A1 VGND VGND VPWR VPWR U$$2625/A1 sky130_fd_sc_hd__buf_4
XFILLER_113_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrepeater1484 U$$3719/A1 VGND VGND VPWR VPWR U$$4402/B1 sky130_fd_sc_hd__buf_4
XFILLER_67_1065 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_956 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater1495 input124/X VGND VGND VPWR VPWR U$$4242/B1 sky130_fd_sc_hd__buf_4
XFILLER_141_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdadda_fa_5_65_1 dadda_fa_5_65_1/A dadda_fa_5_65_1/B dadda_fa_5_65_1/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_66_0/B dadda_fa_7_65_0/A sky130_fd_sc_hd__fa_2
XFILLER_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_1177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xdadda_fa_5_58_0 dadda_fa_5_58_0/A dadda_fa_5_58_0/B dadda_fa_5_58_0/CIN VGND VGND
+ VPWR VPWR dadda_fa_6_59_0/A dadda_fa_6_58_0/CIN sky130_fd_sc_hd__fa_1
XFILLER_140_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
.ends

