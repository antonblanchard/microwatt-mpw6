VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM32_1RW1R
  CLASS BLOCK ;
  FOREIGN RAM32_1RW1R ;
  ORIGIN 0.000 0.000 ;
  SIZE 1173.460 BY 185.440 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 125.160 1173.460 125.760 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 138.760 1173.460 139.360 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 151.680 1173.460 152.280 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 165.280 1173.460 165.880 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 178.200 1173.460 178.800 ;
    END
  END A0[4]
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 2.000 40.080 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 2.000 66.600 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.000 93.120 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 2.000 119.640 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 2.000 146.160 ;
    END
  END A1[4]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.000 13.560 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 2.000 ;
    END
  END Di0[31]
  PIN Di0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 2.000 ;
    END
  END Di0[32]
  PIN Di0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.730 0.000 614.010 2.000 ;
    END
  END Di0[33]
  PIN Di0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 2.000 ;
    END
  END Di0[34]
  PIN Di0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 2.000 ;
    END
  END Di0[35]
  PIN Di0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.470 0.000 668.750 2.000 ;
    END
  END Di0[36]
  PIN Di0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 2.000 ;
    END
  END Di0[37]
  PIN Di0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 2.000 ;
    END
  END Di0[38]
  PIN Di0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 2.000 ;
    END
  END Di0[39]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 2.000 ;
    END
  END Di0[3]
  PIN Di0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 0.000 742.350 2.000 ;
    END
  END Di0[40]
  PIN Di0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 0.000 760.750 2.000 ;
    END
  END Di0[41]
  PIN Di0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 0.000 779.150 2.000 ;
    END
  END Di0[42]
  PIN Di0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 2.000 ;
    END
  END Di0[43]
  PIN Di0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 2.000 ;
    END
  END Di0[44]
  PIN Di0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 0.000 833.890 2.000 ;
    END
  END Di0[45]
  PIN Di0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 0.000 852.290 2.000 ;
    END
  END Di0[46]
  PIN Di0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 2.000 ;
    END
  END Di0[47]
  PIN Di0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 2.000 ;
    END
  END Di0[48]
  PIN Di0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 2.000 ;
    END
  END Di0[49]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 2.000 ;
    END
  END Di0[4]
  PIN Di0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.150 0.000 925.430 2.000 ;
    END
  END Di0[50]
  PIN Di0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 2.000 ;
    END
  END Di0[51]
  PIN Di0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.950 0.000 962.230 2.000 ;
    END
  END Di0[52]
  PIN Di0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 0.000 980.630 2.000 ;
    END
  END Di0[53]
  PIN Di0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 2.000 ;
    END
  END Di0[54]
  PIN Di0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 0.000 1017.430 2.000 ;
    END
  END Di0[55]
  PIN Di0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.550 0.000 1035.830 2.000 ;
    END
  END Di0[56]
  PIN Di0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.490 0.000 1053.770 2.000 ;
    END
  END Di0[57]
  PIN Di0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 0.000 1072.170 2.000 ;
    END
  END Di0[58]
  PIN Di0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.290 0.000 1090.570 2.000 ;
    END
  END Di0[59]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 2.000 ;
    END
  END Di0[5]
  PIN Di0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.690 0.000 1108.970 2.000 ;
    END
  END Di0[60]
  PIN Di0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 2.000 ;
    END
  END Di0[61]
  PIN Di0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.490 0.000 1145.770 2.000 ;
    END
  END Di0[62]
  PIN Di0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 0.000 1164.170 2.000 ;
    END
  END Di0[63]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 183.440 4.510 185.440 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 183.440 96.050 185.440 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 183.440 114.450 185.440 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 183.440 132.850 185.440 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 183.440 150.790 185.440 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 183.440 169.190 185.440 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 183.440 187.590 185.440 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 183.440 205.990 185.440 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 183.440 224.390 185.440 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 183.440 242.790 185.440 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 183.440 261.190 185.440 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 183.440 13.250 185.440 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 183.440 279.130 185.440 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 183.440 288.330 185.440 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 183.440 297.530 185.440 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 183.440 306.730 185.440 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 183.440 315.930 185.440 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 183.440 325.130 185.440 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 183.440 334.330 185.440 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 183.440 343.530 185.440 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 183.440 352.730 185.440 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 183.440 361.930 185.440 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 183.440 22.450 185.440 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 183.440 371.130 185.440 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 183.440 380.330 185.440 ;
    END
  END Do0[31]
  PIN Do0[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 183.440 389.530 185.440 ;
    END
  END Do0[32]
  PIN Do0[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 183.440 398.270 185.440 ;
    END
  END Do0[33]
  PIN Do0[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 183.440 407.470 185.440 ;
    END
  END Do0[34]
  PIN Do0[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 183.440 416.670 185.440 ;
    END
  END Do0[35]
  PIN Do0[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 183.440 425.870 185.440 ;
    END
  END Do0[36]
  PIN Do0[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 183.440 435.070 185.440 ;
    END
  END Do0[37]
  PIN Do0[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 183.440 444.270 185.440 ;
    END
  END Do0[38]
  PIN Do0[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 183.440 453.470 185.440 ;
    END
  END Do0[39]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 183.440 31.650 185.440 ;
    END
  END Do0[3]
  PIN Do0[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 183.440 462.670 185.440 ;
    END
  END Do0[40]
  PIN Do0[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 183.440 471.870 185.440 ;
    END
  END Do0[41]
  PIN Do0[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 183.440 481.070 185.440 ;
    END
  END Do0[42]
  PIN Do0[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 183.440 490.270 185.440 ;
    END
  END Do0[43]
  PIN Do0[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 183.440 499.470 185.440 ;
    END
  END Do0[44]
  PIN Do0[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 183.440 508.670 185.440 ;
    END
  END Do0[45]
  PIN Do0[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 183.440 517.870 185.440 ;
    END
  END Do0[46]
  PIN Do0[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 183.440 526.610 185.440 ;
    END
  END Do0[47]
  PIN Do0[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 183.440 535.810 185.440 ;
    END
  END Do0[48]
  PIN Do0[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 183.440 545.010 185.440 ;
    END
  END Do0[49]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 183.440 40.850 185.440 ;
    END
  END Do0[4]
  PIN Do0[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 183.440 554.210 185.440 ;
    END
  END Do0[50]
  PIN Do0[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 183.440 563.410 185.440 ;
    END
  END Do0[51]
  PIN Do0[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 183.440 572.610 185.440 ;
    END
  END Do0[52]
  PIN Do0[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 183.440 581.810 185.440 ;
    END
  END Do0[53]
  PIN Do0[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 183.440 591.010 185.440 ;
    END
  END Do0[54]
  PIN Do0[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 183.440 600.210 185.440 ;
    END
  END Do0[55]
  PIN Do0[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 183.440 609.410 185.440 ;
    END
  END Do0[56]
  PIN Do0[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 183.440 618.610 185.440 ;
    END
  END Do0[57]
  PIN Do0[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 183.440 627.810 185.440 ;
    END
  END Do0[58]
  PIN Do0[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 183.440 637.010 185.440 ;
    END
  END Do0[59]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 183.440 50.050 185.440 ;
    END
  END Do0[5]
  PIN Do0[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 183.440 646.210 185.440 ;
    END
  END Do0[60]
  PIN Do0[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 183.440 655.410 185.440 ;
    END
  END Do0[61]
  PIN Do0[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 183.440 664.150 185.440 ;
    END
  END Do0[62]
  PIN Do0[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 183.440 673.350 185.440 ;
    END
  END Do0[63]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 183.440 59.250 185.440 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 183.440 68.450 185.440 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 183.440 77.650 185.440 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 183.440 86.850 185.440 ;
    END
  END Do0[9]
  PIN Do1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 183.440 105.250 185.440 ;
    END
  END Do1[0]
  PIN Do1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 183.440 682.550 185.440 ;
    END
  END Do1[10]
  PIN Do1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 183.440 691.750 185.440 ;
    END
  END Do1[11]
  PIN Do1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 183.440 700.950 185.440 ;
    END
  END Do1[12]
  PIN Do1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.870 183.440 710.150 185.440 ;
    END
  END Do1[13]
  PIN Do1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 183.440 719.350 185.440 ;
    END
  END Do1[14]
  PIN Do1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 183.440 728.550 185.440 ;
    END
  END Do1[15]
  PIN Do1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 183.440 737.750 185.440 ;
    END
  END Do1[16]
  PIN Do1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 183.440 746.950 185.440 ;
    END
  END Do1[17]
  PIN Do1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 183.440 756.150 185.440 ;
    END
  END Do1[18]
  PIN Do1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.070 183.440 765.350 185.440 ;
    END
  END Do1[19]
  PIN Do1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 183.440 123.650 185.440 ;
    END
  END Do1[1]
  PIN Do1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.270 183.440 774.550 185.440 ;
    END
  END Do1[20]
  PIN Do1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 183.440 783.750 185.440 ;
    END
  END Do1[21]
  PIN Do1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 183.440 792.490 185.440 ;
    END
  END Do1[22]
  PIN Do1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 183.440 801.690 185.440 ;
    END
  END Do1[23]
  PIN Do1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 183.440 810.890 185.440 ;
    END
  END Do1[24]
  PIN Do1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 183.440 820.090 185.440 ;
    END
  END Do1[25]
  PIN Do1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 183.440 829.290 185.440 ;
    END
  END Do1[26]
  PIN Do1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 183.440 838.490 185.440 ;
    END
  END Do1[27]
  PIN Do1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 183.440 847.690 185.440 ;
    END
  END Do1[28]
  PIN Do1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 183.440 856.890 185.440 ;
    END
  END Do1[29]
  PIN Do1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 183.440 141.590 185.440 ;
    END
  END Do1[2]
  PIN Do1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 183.440 866.090 185.440 ;
    END
  END Do1[30]
  PIN Do1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 183.440 875.290 185.440 ;
    END
  END Do1[31]
  PIN Do1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.210 183.440 884.490 185.440 ;
    END
  END Do1[32]
  PIN Do1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 183.440 893.690 185.440 ;
    END
  END Do1[33]
  PIN Do1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 183.440 902.890 185.440 ;
    END
  END Do1[34]
  PIN Do1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 183.440 912.090 185.440 ;
    END
  END Do1[35]
  PIN Do1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 183.440 920.830 185.440 ;
    END
  END Do1[36]
  PIN Do1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 183.440 930.030 185.440 ;
    END
  END Do1[37]
  PIN Do1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.950 183.440 939.230 185.440 ;
    END
  END Do1[38]
  PIN Do1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 183.440 948.430 185.440 ;
    END
  END Do1[39]
  PIN Do1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 183.440 159.990 185.440 ;
    END
  END Do1[3]
  PIN Do1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 183.440 957.630 185.440 ;
    END
  END Do1[40]
  PIN Do1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 183.440 966.830 185.440 ;
    END
  END Do1[41]
  PIN Do1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 183.440 976.030 185.440 ;
    END
  END Do1[42]
  PIN Do1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 183.440 985.230 185.440 ;
    END
  END Do1[43]
  PIN Do1[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.150 183.440 994.430 185.440 ;
    END
  END Do1[44]
  PIN Do1[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.350 183.440 1003.630 185.440 ;
    END
  END Do1[45]
  PIN Do1[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.550 183.440 1012.830 185.440 ;
    END
  END Do1[46]
  PIN Do1[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.750 183.440 1022.030 185.440 ;
    END
  END Do1[47]
  PIN Do1[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 183.440 1031.230 185.440 ;
    END
  END Do1[48]
  PIN Do1[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 183.440 1040.430 185.440 ;
    END
  END Do1[49]
  PIN Do1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 183.440 178.390 185.440 ;
    END
  END Do1[4]
  PIN Do1[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.890 183.440 1049.170 185.440 ;
    END
  END Do1[50]
  PIN Do1[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 183.440 1058.370 185.440 ;
    END
  END Do1[51]
  PIN Do1[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.290 183.440 1067.570 185.440 ;
    END
  END Do1[52]
  PIN Do1[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 183.440 1076.770 185.440 ;
    END
  END Do1[53]
  PIN Do1[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.690 183.440 1085.970 185.440 ;
    END
  END Do1[54]
  PIN Do1[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 183.440 1095.170 185.440 ;
    END
  END Do1[55]
  PIN Do1[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 183.440 1104.370 185.440 ;
    END
  END Do1[56]
  PIN Do1[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.290 183.440 1113.570 185.440 ;
    END
  END Do1[57]
  PIN Do1[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.490 183.440 1122.770 185.440 ;
    END
  END Do1[58]
  PIN Do1[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.690 183.440 1131.970 185.440 ;
    END
  END Do1[59]
  PIN Do1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 183.440 196.790 185.440 ;
    END
  END Do1[5]
  PIN Do1[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.890 183.440 1141.170 185.440 ;
    END
  END Do1[60]
  PIN Do1[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 183.440 1150.370 185.440 ;
    END
  END Do1[61]
  PIN Do1[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 183.440 1159.570 185.440 ;
    END
  END Do1[62]
  PIN Do1[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.490 183.440 1168.770 185.440 ;
    END
  END Do1[63]
  PIN Do1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 183.440 215.190 185.440 ;
    END
  END Do1[6]
  PIN Do1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 183.440 233.590 185.440 ;
    END
  END Do1[7]
  PIN Do1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 183.440 251.990 185.440 ;
    END
  END Do1[8]
  PIN Do1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 183.440 269.930 185.440 ;
    END
  END Do1[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 6.160 1173.460 6.760 ;
    END
  END EN0
  PIN EN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 2.000 172.680 ;
    END
  END EN1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.210 2.480 99.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.210 2.480 279.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 456.210 2.480 459.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.210 2.480 639.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 816.210 2.480 819.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 996.210 2.480 999.310 182.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 6.210 2.480 9.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 186.210 2.480 189.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 366.210 2.480 369.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 546.210 2.480 549.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 726.210 2.480 729.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 906.210 2.480 909.310 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1086.210 2.480 1089.310 182.480 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 19.080 1173.460 19.680 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 32.680 1173.460 33.280 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 45.600 1173.460 46.200 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 59.200 1173.460 59.800 ;
    END
  END WE0[3]
  PIN WE0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 72.120 1173.460 72.720 ;
    END
  END WE0[4]
  PIN WE0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 85.720 1173.460 86.320 ;
    END
  END WE0[5]
  PIN WE0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 98.640 1173.460 99.240 ;
    END
  END WE0[6]
  PIN WE0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1171.460 112.240 1173.460 112.840 ;
    END
  END WE0[7]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 1170.700 98.005 ;
      LAYER met1 ;
        RECT 0.990 0.380 1170.700 183.560 ;
      LAYER met2 ;
        RECT 1.020 183.160 3.950 184.010 ;
        RECT 4.790 183.160 12.690 184.010 ;
        RECT 13.530 183.160 21.890 184.010 ;
        RECT 22.730 183.160 31.090 184.010 ;
        RECT 31.930 183.160 40.290 184.010 ;
        RECT 41.130 183.160 49.490 184.010 ;
        RECT 50.330 183.160 58.690 184.010 ;
        RECT 59.530 183.160 67.890 184.010 ;
        RECT 68.730 183.160 77.090 184.010 ;
        RECT 77.930 183.160 86.290 184.010 ;
        RECT 87.130 183.160 95.490 184.010 ;
        RECT 96.330 183.160 104.690 184.010 ;
        RECT 105.530 183.160 113.890 184.010 ;
        RECT 114.730 183.160 123.090 184.010 ;
        RECT 123.930 183.160 132.290 184.010 ;
        RECT 133.130 183.160 141.030 184.010 ;
        RECT 141.870 183.160 150.230 184.010 ;
        RECT 151.070 183.160 159.430 184.010 ;
        RECT 160.270 183.160 168.630 184.010 ;
        RECT 169.470 183.160 177.830 184.010 ;
        RECT 178.670 183.160 187.030 184.010 ;
        RECT 187.870 183.160 196.230 184.010 ;
        RECT 197.070 183.160 205.430 184.010 ;
        RECT 206.270 183.160 214.630 184.010 ;
        RECT 215.470 183.160 223.830 184.010 ;
        RECT 224.670 183.160 233.030 184.010 ;
        RECT 233.870 183.160 242.230 184.010 ;
        RECT 243.070 183.160 251.430 184.010 ;
        RECT 252.270 183.160 260.630 184.010 ;
        RECT 261.470 183.160 269.370 184.010 ;
        RECT 270.210 183.160 278.570 184.010 ;
        RECT 279.410 183.160 287.770 184.010 ;
        RECT 288.610 183.160 296.970 184.010 ;
        RECT 297.810 183.160 306.170 184.010 ;
        RECT 307.010 183.160 315.370 184.010 ;
        RECT 316.210 183.160 324.570 184.010 ;
        RECT 325.410 183.160 333.770 184.010 ;
        RECT 334.610 183.160 342.970 184.010 ;
        RECT 343.810 183.160 352.170 184.010 ;
        RECT 353.010 183.160 361.370 184.010 ;
        RECT 362.210 183.160 370.570 184.010 ;
        RECT 371.410 183.160 379.770 184.010 ;
        RECT 380.610 183.160 388.970 184.010 ;
        RECT 389.810 183.160 397.710 184.010 ;
        RECT 398.550 183.160 406.910 184.010 ;
        RECT 407.750 183.160 416.110 184.010 ;
        RECT 416.950 183.160 425.310 184.010 ;
        RECT 426.150 183.160 434.510 184.010 ;
        RECT 435.350 183.160 443.710 184.010 ;
        RECT 444.550 183.160 452.910 184.010 ;
        RECT 453.750 183.160 462.110 184.010 ;
        RECT 462.950 183.160 471.310 184.010 ;
        RECT 472.150 183.160 480.510 184.010 ;
        RECT 481.350 183.160 489.710 184.010 ;
        RECT 490.550 183.160 498.910 184.010 ;
        RECT 499.750 183.160 508.110 184.010 ;
        RECT 508.950 183.160 517.310 184.010 ;
        RECT 518.150 183.160 526.050 184.010 ;
        RECT 526.890 183.160 535.250 184.010 ;
        RECT 536.090 183.160 544.450 184.010 ;
        RECT 545.290 183.160 553.650 184.010 ;
        RECT 554.490 183.160 562.850 184.010 ;
        RECT 563.690 183.160 572.050 184.010 ;
        RECT 572.890 183.160 581.250 184.010 ;
        RECT 582.090 183.160 590.450 184.010 ;
        RECT 591.290 183.160 599.650 184.010 ;
        RECT 600.490 183.160 608.850 184.010 ;
        RECT 609.690 183.160 618.050 184.010 ;
        RECT 618.890 183.160 627.250 184.010 ;
        RECT 628.090 183.160 636.450 184.010 ;
        RECT 637.290 183.160 645.650 184.010 ;
        RECT 646.490 183.160 654.850 184.010 ;
        RECT 655.690 183.160 663.590 184.010 ;
        RECT 664.430 183.160 672.790 184.010 ;
        RECT 673.630 183.160 681.990 184.010 ;
        RECT 682.830 183.160 691.190 184.010 ;
        RECT 692.030 183.160 700.390 184.010 ;
        RECT 701.230 183.160 709.590 184.010 ;
        RECT 710.430 183.160 718.790 184.010 ;
        RECT 719.630 183.160 727.990 184.010 ;
        RECT 728.830 183.160 737.190 184.010 ;
        RECT 738.030 183.160 746.390 184.010 ;
        RECT 747.230 183.160 755.590 184.010 ;
        RECT 756.430 183.160 764.790 184.010 ;
        RECT 765.630 183.160 773.990 184.010 ;
        RECT 774.830 183.160 783.190 184.010 ;
        RECT 784.030 183.160 791.930 184.010 ;
        RECT 792.770 183.160 801.130 184.010 ;
        RECT 801.970 183.160 810.330 184.010 ;
        RECT 811.170 183.160 819.530 184.010 ;
        RECT 820.370 183.160 828.730 184.010 ;
        RECT 829.570 183.160 837.930 184.010 ;
        RECT 838.770 183.160 847.130 184.010 ;
        RECT 847.970 183.160 856.330 184.010 ;
        RECT 857.170 183.160 865.530 184.010 ;
        RECT 866.370 183.160 874.730 184.010 ;
        RECT 875.570 183.160 883.930 184.010 ;
        RECT 884.770 183.160 893.130 184.010 ;
        RECT 893.970 183.160 902.330 184.010 ;
        RECT 903.170 183.160 911.530 184.010 ;
        RECT 912.370 183.160 920.270 184.010 ;
        RECT 921.110 183.160 929.470 184.010 ;
        RECT 930.310 183.160 938.670 184.010 ;
        RECT 939.510 183.160 947.870 184.010 ;
        RECT 948.710 183.160 957.070 184.010 ;
        RECT 957.910 183.160 966.270 184.010 ;
        RECT 967.110 183.160 975.470 184.010 ;
        RECT 976.310 183.160 984.670 184.010 ;
        RECT 985.510 183.160 993.870 184.010 ;
        RECT 994.710 183.160 1003.070 184.010 ;
        RECT 1003.910 183.160 1012.270 184.010 ;
        RECT 1013.110 183.160 1021.470 184.010 ;
        RECT 1022.310 183.160 1030.670 184.010 ;
        RECT 1031.510 183.160 1039.870 184.010 ;
        RECT 1040.710 183.160 1048.610 184.010 ;
        RECT 1049.450 183.160 1057.810 184.010 ;
        RECT 1058.650 183.160 1067.010 184.010 ;
        RECT 1067.850 183.160 1076.210 184.010 ;
        RECT 1077.050 183.160 1085.410 184.010 ;
        RECT 1086.250 183.160 1094.610 184.010 ;
        RECT 1095.450 183.160 1103.810 184.010 ;
        RECT 1104.650 183.160 1113.010 184.010 ;
        RECT 1113.850 183.160 1122.210 184.010 ;
        RECT 1123.050 183.160 1131.410 184.010 ;
        RECT 1132.250 183.160 1140.610 184.010 ;
        RECT 1141.450 183.160 1149.810 184.010 ;
        RECT 1150.650 183.160 1159.010 184.010 ;
        RECT 1159.850 183.160 1168.210 184.010 ;
        RECT 1169.050 183.160 1169.680 184.010 ;
        RECT 1.020 2.280 1169.680 183.160 ;
        RECT 1.020 0.155 8.550 2.280 ;
        RECT 9.390 0.155 26.490 2.280 ;
        RECT 27.330 0.155 44.890 2.280 ;
        RECT 45.730 0.155 63.290 2.280 ;
        RECT 64.130 0.155 81.690 2.280 ;
        RECT 82.530 0.155 100.090 2.280 ;
        RECT 100.930 0.155 118.490 2.280 ;
        RECT 119.330 0.155 136.890 2.280 ;
        RECT 137.730 0.155 154.830 2.280 ;
        RECT 155.670 0.155 173.230 2.280 ;
        RECT 174.070 0.155 191.630 2.280 ;
        RECT 192.470 0.155 210.030 2.280 ;
        RECT 210.870 0.155 228.430 2.280 ;
        RECT 229.270 0.155 246.830 2.280 ;
        RECT 247.670 0.155 265.230 2.280 ;
        RECT 266.070 0.155 283.170 2.280 ;
        RECT 284.010 0.155 301.570 2.280 ;
        RECT 302.410 0.155 319.970 2.280 ;
        RECT 320.810 0.155 338.370 2.280 ;
        RECT 339.210 0.155 356.770 2.280 ;
        RECT 357.610 0.155 375.170 2.280 ;
        RECT 376.010 0.155 393.570 2.280 ;
        RECT 394.410 0.155 411.510 2.280 ;
        RECT 412.350 0.155 429.910 2.280 ;
        RECT 430.750 0.155 448.310 2.280 ;
        RECT 449.150 0.155 466.710 2.280 ;
        RECT 467.550 0.155 485.110 2.280 ;
        RECT 485.950 0.155 503.510 2.280 ;
        RECT 504.350 0.155 521.910 2.280 ;
        RECT 522.750 0.155 539.850 2.280 ;
        RECT 540.690 0.155 558.250 2.280 ;
        RECT 559.090 0.155 576.650 2.280 ;
        RECT 577.490 0.155 595.050 2.280 ;
        RECT 595.890 0.155 613.450 2.280 ;
        RECT 614.290 0.155 631.850 2.280 ;
        RECT 632.690 0.155 650.250 2.280 ;
        RECT 651.090 0.155 668.190 2.280 ;
        RECT 669.030 0.155 686.590 2.280 ;
        RECT 687.430 0.155 704.990 2.280 ;
        RECT 705.830 0.155 723.390 2.280 ;
        RECT 724.230 0.155 741.790 2.280 ;
        RECT 742.630 0.155 760.190 2.280 ;
        RECT 761.030 0.155 778.590 2.280 ;
        RECT 779.430 0.155 796.530 2.280 ;
        RECT 797.370 0.155 814.930 2.280 ;
        RECT 815.770 0.155 833.330 2.280 ;
        RECT 834.170 0.155 851.730 2.280 ;
        RECT 852.570 0.155 870.130 2.280 ;
        RECT 870.970 0.155 888.530 2.280 ;
        RECT 889.370 0.155 906.930 2.280 ;
        RECT 907.770 0.155 924.870 2.280 ;
        RECT 925.710 0.155 943.270 2.280 ;
        RECT 944.110 0.155 961.670 2.280 ;
        RECT 962.510 0.155 980.070 2.280 ;
        RECT 980.910 0.155 998.470 2.280 ;
        RECT 999.310 0.155 1016.870 2.280 ;
        RECT 1017.710 0.155 1035.270 2.280 ;
        RECT 1036.110 0.155 1053.210 2.280 ;
        RECT 1054.050 0.155 1071.610 2.280 ;
        RECT 1072.450 0.155 1090.010 2.280 ;
        RECT 1090.850 0.155 1108.410 2.280 ;
        RECT 1109.250 0.155 1126.810 2.280 ;
        RECT 1127.650 0.155 1145.210 2.280 ;
        RECT 1146.050 0.155 1163.610 2.280 ;
        RECT 1164.450 0.155 1169.680 2.280 ;
      LAYER met3 ;
        RECT 1.905 179.200 1171.460 182.405 ;
        RECT 1.905 177.800 1171.060 179.200 ;
        RECT 1.905 173.080 1171.460 177.800 ;
        RECT 2.400 171.680 1171.460 173.080 ;
        RECT 1.905 166.280 1171.460 171.680 ;
        RECT 1.905 164.880 1171.060 166.280 ;
        RECT 1.905 152.680 1171.460 164.880 ;
        RECT 1.905 151.280 1171.060 152.680 ;
        RECT 1.905 146.560 1171.460 151.280 ;
        RECT 2.400 145.160 1171.460 146.560 ;
        RECT 1.905 139.760 1171.460 145.160 ;
        RECT 1.905 138.360 1171.060 139.760 ;
        RECT 1.905 126.160 1171.460 138.360 ;
        RECT 1.905 124.760 1171.060 126.160 ;
        RECT 1.905 120.040 1171.460 124.760 ;
        RECT 2.400 118.640 1171.460 120.040 ;
        RECT 1.905 113.240 1171.460 118.640 ;
        RECT 1.905 111.840 1171.060 113.240 ;
        RECT 1.905 99.640 1171.460 111.840 ;
        RECT 1.905 98.240 1171.060 99.640 ;
        RECT 1.905 93.520 1171.460 98.240 ;
        RECT 2.400 92.120 1171.460 93.520 ;
        RECT 1.905 86.720 1171.460 92.120 ;
        RECT 1.905 85.320 1171.060 86.720 ;
        RECT 1.905 73.120 1171.460 85.320 ;
        RECT 1.905 71.720 1171.060 73.120 ;
        RECT 1.905 67.000 1171.460 71.720 ;
        RECT 2.400 65.600 1171.460 67.000 ;
        RECT 1.905 60.200 1171.460 65.600 ;
        RECT 1.905 58.800 1171.060 60.200 ;
        RECT 1.905 46.600 1171.460 58.800 ;
        RECT 1.905 45.200 1171.060 46.600 ;
        RECT 1.905 40.480 1171.460 45.200 ;
        RECT 2.400 39.080 1171.460 40.480 ;
        RECT 1.905 33.680 1171.460 39.080 ;
        RECT 1.905 32.280 1171.060 33.680 ;
        RECT 1.905 20.080 1171.460 32.280 ;
        RECT 1.905 18.680 1171.060 20.080 ;
        RECT 1.905 13.960 1171.460 18.680 ;
        RECT 2.400 12.560 1171.460 13.960 ;
        RECT 1.905 7.160 1171.460 12.560 ;
        RECT 1.905 5.760 1171.060 7.160 ;
        RECT 1.905 0.175 1171.460 5.760 ;
      LAYER met4 ;
        RECT 4.895 2.080 5.810 177.985 ;
        RECT 9.710 2.080 95.810 177.985 ;
        RECT 99.710 2.080 185.810 177.985 ;
        RECT 189.710 2.080 275.810 177.985 ;
        RECT 279.710 2.080 365.810 177.985 ;
        RECT 369.710 2.080 455.810 177.985 ;
        RECT 459.710 2.080 545.810 177.985 ;
        RECT 549.710 2.080 635.810 177.985 ;
        RECT 639.710 2.080 725.810 177.985 ;
        RECT 729.710 2.080 815.810 177.985 ;
        RECT 819.710 2.080 905.810 177.985 ;
        RECT 909.710 2.080 995.810 177.985 ;
        RECT 999.710 2.080 1077.945 177.985 ;
        RECT 4.895 0.855 1077.945 2.080 ;
  END
END RAM32_1RW1R
END LIBRARY

